magic
tech scmos
magscale 1 2
timestamp 1745250350
<< metal1 >>
rect 680 2006 686 2014
rect 694 2006 700 2014
rect 708 2006 714 2014
rect 722 2006 728 2014
rect 1117 1917 1139 1923
rect 1236 1916 1244 1924
rect 957 1897 972 1903
rect 1181 1897 1235 1903
rect 1268 1897 1283 1903
rect 1758 1897 1843 1903
rect 1892 1897 1907 1903
rect 1053 1877 1080 1883
rect 1917 1877 1932 1883
rect 781 1857 812 1863
rect 2349 1857 2380 1863
rect 1688 1806 1694 1814
rect 1702 1806 1708 1814
rect 1716 1806 1722 1814
rect 1730 1806 1736 1814
rect 72 1776 76 1784
rect 2084 1776 2088 1784
rect 740 1757 764 1763
rect 804 1757 819 1763
rect 1108 1757 1139 1763
rect 2317 1757 2332 1763
rect 446 1737 483 1743
rect 573 1723 579 1743
rect 637 1737 700 1743
rect 900 1737 915 1743
rect 1069 1737 1091 1743
rect 1629 1737 1676 1743
rect 2157 1743 2163 1756
rect 2014 1737 2051 1743
rect 2141 1737 2163 1743
rect 2365 1743 2371 1763
rect 2292 1737 2307 1743
rect 2365 1737 2403 1743
rect 468 1717 520 1723
rect 573 1717 611 1723
rect 845 1717 883 1723
rect 1037 1717 1068 1723
rect 1588 1717 1619 1723
rect 2189 1717 2227 1723
rect 2269 1717 2284 1723
rect 621 1697 643 1703
rect 893 1697 908 1703
rect 1124 1697 1139 1703
rect 836 1636 838 1644
rect 680 1606 686 1614
rect 694 1606 700 1614
rect 708 1606 714 1614
rect 722 1606 728 1614
rect 2381 1537 2396 1543
rect 852 1516 856 1524
rect 1284 1477 1299 1483
rect 1837 1477 1852 1483
rect 2212 1477 2227 1483
rect 685 1457 716 1463
rect 2237 1457 2275 1463
rect 1780 1436 1784 1444
rect 1688 1406 1694 1414
rect 1702 1406 1708 1414
rect 1716 1406 1722 1414
rect 1730 1406 1736 1414
rect 452 1376 456 1384
rect 936 1376 940 1384
rect 1976 1376 1980 1384
rect 724 1357 755 1363
rect 765 1357 780 1363
rect 1229 1357 1260 1363
rect 1821 1357 1843 1363
rect 509 1337 547 1343
rect 797 1337 828 1343
rect 1341 1337 1363 1343
rect 1805 1317 1820 1323
rect 636 1312 644 1316
rect 621 1297 643 1303
rect 1860 1297 1875 1303
rect 588 1292 596 1296
rect 68 1277 83 1283
rect 680 1206 686 1214
rect 694 1206 700 1214
rect 708 1206 714 1214
rect 722 1206 728 1214
rect 1133 1137 1164 1143
rect 1820 1132 1828 1136
rect 45 1097 82 1103
rect 733 1097 748 1103
rect 877 1097 892 1103
rect 1805 1097 1843 1103
rect 2190 1097 2227 1103
rect 1668 1077 1731 1083
rect 1780 1077 1795 1083
rect 589 1057 620 1063
rect 1748 1057 1779 1063
rect 452 1036 456 1044
rect 941 1037 956 1043
rect 1172 1037 1187 1043
rect 1688 1006 1694 1014
rect 1702 1006 1708 1014
rect 1716 1006 1722 1014
rect 1730 1006 1736 1014
rect 788 977 803 983
rect 1210 976 1212 984
rect 1290 976 1292 984
rect 1565 957 1580 963
rect 2301 957 2316 963
rect 468 937 483 943
rect 1005 937 1052 943
rect 1069 937 1100 943
rect 1140 937 1155 943
rect 1165 937 1196 943
rect 1229 937 1244 943
rect 1437 937 1484 943
rect 1805 937 1827 943
rect 653 917 723 923
rect 1236 917 1251 923
rect 1309 917 1331 923
rect 1428 917 1507 923
rect 1773 917 1788 923
rect 1853 917 1868 923
rect 2324 917 2339 923
rect 1869 897 1891 903
rect 1196 884 1204 888
rect 1604 877 1619 883
rect 1645 877 1724 883
rect 1645 857 1651 877
rect 2365 877 2396 883
rect 680 806 686 814
rect 694 806 700 814
rect 708 806 714 814
rect 722 806 728 814
rect 2301 737 2316 743
rect 45 697 82 703
rect 1229 697 1276 703
rect 1261 677 1298 683
rect 1768 676 1772 684
rect 1949 677 1964 683
rect 2365 677 2396 683
rect 1837 657 1852 663
rect 1688 606 1694 614
rect 1702 606 1708 614
rect 1716 606 1722 614
rect 1730 606 1736 614
rect 413 557 444 563
rect 541 557 572 563
rect 388 537 403 543
rect 468 537 483 543
rect 637 543 643 563
rect 989 557 1004 563
rect 637 537 675 543
rect 724 537 771 543
rect 61 523 67 536
rect 1037 543 1043 556
rect 916 537 931 543
rect 1037 537 1059 543
rect 1197 537 1235 543
rect 1796 537 1811 543
rect 45 517 67 523
rect 157 517 179 523
rect 372 517 387 523
rect 685 517 748 523
rect 893 517 924 523
rect 1021 517 1052 523
rect 1821 517 1859 523
rect 509 497 531 503
rect 957 497 972 503
rect 1101 497 1123 503
rect 1924 496 1932 504
rect 525 477 540 483
rect 1252 477 1283 483
rect 680 406 686 414
rect 694 406 700 414
rect 708 406 714 414
rect 722 406 728 414
rect 2077 317 2099 323
rect 756 297 856 303
rect 909 297 924 303
rect 734 277 812 283
rect 909 277 915 297
rect 941 297 979 303
rect 1116 292 1124 296
rect 1053 277 1068 283
rect 1085 277 1123 283
rect 1197 277 1235 283
rect 1005 257 1036 263
rect 1229 257 1235 277
rect 1965 277 1980 283
rect 1788 264 1796 268
rect 1245 257 1276 263
rect 2004 257 2035 263
rect 1908 236 1912 244
rect 1688 206 1694 214
rect 1702 206 1708 214
rect 1716 206 1722 214
rect 1730 206 1736 214
rect 1320 176 1324 184
rect 420 117 451 123
rect 1060 117 1075 123
rect 1085 117 1107 123
rect 1357 123 1363 136
rect 1357 117 1379 123
rect 1516 117 1555 123
rect 1516 116 1524 117
rect 680 6 686 14
rect 694 6 700 14
rect 708 6 714 14
rect 722 6 728 14
<< m2contact >>
rect 686 2006 694 2014
rect 700 2006 708 2014
rect 714 2006 722 2014
rect 316 1976 324 1984
rect 396 1976 404 1984
rect 444 1976 452 1984
rect 492 1976 500 1984
rect 860 1976 868 1984
rect 1308 1976 1316 1984
rect 1356 1976 1364 1984
rect 1468 1976 1476 1984
rect 1868 1976 1876 1984
rect 2012 1976 2020 1984
rect 2060 1976 2068 1984
rect 1084 1936 1092 1944
rect 316 1916 324 1924
rect 492 1916 500 1924
rect 972 1916 980 1924
rect 1020 1916 1028 1924
rect 1196 1916 1204 1924
rect 1228 1916 1236 1924
rect 1260 1916 1268 1924
rect 1468 1916 1476 1924
rect 1884 1916 1892 1924
rect 1932 1916 1940 1924
rect 2060 1916 2068 1924
rect 316 1896 324 1904
rect 364 1896 372 1904
rect 412 1896 420 1904
rect 492 1896 500 1904
rect 892 1896 900 1904
rect 924 1896 932 1904
rect 972 1896 980 1904
rect 1100 1896 1108 1904
rect 1260 1896 1268 1904
rect 1324 1896 1332 1904
rect 1388 1896 1396 1904
rect 1420 1896 1428 1904
rect 1468 1896 1476 1904
rect 1884 1896 1892 1904
rect 1980 1896 1988 1904
rect 2060 1896 2068 1904
rect 220 1876 228 1884
rect 588 1876 596 1884
rect 908 1876 916 1884
rect 1004 1876 1012 1884
rect 1164 1876 1172 1884
rect 1212 1876 1220 1884
rect 1404 1876 1412 1884
rect 1564 1876 1572 1884
rect 1932 1876 1940 1884
rect 1964 1876 1972 1884
rect 2156 1876 2164 1884
rect 188 1856 196 1864
rect 620 1856 628 1864
rect 812 1856 820 1864
rect 1148 1856 1156 1864
rect 1372 1856 1380 1864
rect 1596 1856 1604 1864
rect 2188 1856 2196 1864
rect 2380 1856 2388 1864
rect 28 1836 36 1844
rect 972 1836 980 1844
rect 1020 1836 1028 1844
rect 1756 1836 1764 1844
rect 1932 1836 1940 1844
rect 1694 1806 1702 1814
rect 1708 1806 1716 1814
rect 1722 1806 1730 1814
rect 76 1776 84 1784
rect 444 1776 452 1784
rect 780 1776 788 1784
rect 956 1776 964 1784
rect 1084 1776 1092 1784
rect 1500 1776 1508 1784
rect 1516 1776 1524 1784
rect 2012 1776 2020 1784
rect 2076 1776 2084 1784
rect 2172 1776 2180 1784
rect 284 1756 292 1764
rect 652 1756 660 1764
rect 764 1756 772 1764
rect 796 1756 804 1764
rect 1100 1756 1108 1764
rect 1292 1756 1300 1764
rect 1532 1756 1540 1764
rect 1580 1756 1588 1764
rect 1852 1756 1860 1764
rect 2156 1756 2164 1764
rect 2204 1756 2212 1764
rect 2332 1756 2340 1764
rect 2348 1756 2356 1764
rect 12 1736 20 1744
rect 108 1736 116 1744
rect 252 1736 260 1744
rect 364 1716 372 1724
rect 460 1716 468 1724
rect 588 1736 596 1744
rect 700 1736 708 1744
rect 716 1736 724 1744
rect 860 1736 868 1744
rect 892 1736 900 1744
rect 972 1736 980 1744
rect 1324 1736 1332 1744
rect 1676 1736 1684 1744
rect 1820 1736 1828 1744
rect 2252 1736 2260 1744
rect 2284 1736 2292 1744
rect 2380 1756 2388 1764
rect 764 1716 772 1724
rect 924 1716 932 1724
rect 1068 1716 1076 1724
rect 1212 1716 1220 1724
rect 1436 1716 1444 1724
rect 1468 1716 1476 1724
rect 1548 1716 1556 1724
rect 1580 1716 1588 1724
rect 1724 1716 1732 1724
rect 1932 1716 1940 1724
rect 2236 1716 2244 1724
rect 2284 1716 2292 1724
rect 2332 1716 2340 1724
rect 156 1696 164 1704
rect 748 1696 756 1704
rect 908 1696 916 1704
rect 1116 1696 1124 1704
rect 1388 1700 1396 1708
rect 1596 1696 1604 1704
rect 1756 1700 1764 1708
rect 2284 1696 2292 1704
rect 1388 1654 1396 1662
rect 1756 1654 1764 1662
rect 156 1636 164 1644
rect 828 1636 836 1644
rect 1548 1636 1556 1644
rect 686 1606 694 1614
rect 700 1606 708 1614
rect 714 1606 722 1614
rect 316 1576 324 1584
rect 396 1576 404 1584
rect 764 1576 772 1584
rect 1228 1576 1236 1584
rect 1356 1576 1364 1584
rect 1644 1576 1652 1584
rect 1868 1576 1876 1584
rect 2156 1576 2164 1584
rect 2396 1536 2404 1544
rect 316 1516 324 1524
rect 396 1516 404 1524
rect 844 1516 852 1524
rect 1228 1516 1236 1524
rect 1644 1516 1652 1524
rect 2156 1516 2164 1524
rect 316 1496 324 1504
rect 396 1496 404 1504
rect 796 1496 804 1504
rect 938 1496 946 1504
rect 1212 1496 1220 1504
rect 1228 1496 1236 1504
rect 1324 1496 1332 1504
rect 1436 1496 1444 1504
rect 1948 1496 1956 1504
rect 2204 1496 2212 1504
rect 2252 1496 2260 1504
rect 2300 1496 2308 1504
rect 2348 1496 2356 1504
rect 220 1476 228 1484
rect 492 1476 500 1484
rect 812 1476 820 1484
rect 908 1476 916 1484
rect 1132 1476 1140 1484
rect 1276 1476 1284 1484
rect 1548 1476 1556 1484
rect 1740 1476 1748 1484
rect 1852 1476 1860 1484
rect 2060 1476 2068 1484
rect 2204 1476 2212 1484
rect 2332 1476 2340 1484
rect 188 1456 196 1464
rect 524 1456 532 1464
rect 716 1456 724 1464
rect 1100 1456 1108 1464
rect 1516 1456 1524 1464
rect 2028 1456 2036 1464
rect 2284 1456 2292 1464
rect 28 1436 36 1444
rect 1356 1436 1364 1444
rect 1772 1436 1780 1444
rect 1694 1406 1702 1414
rect 1708 1406 1716 1414
rect 1722 1406 1730 1414
rect 444 1376 452 1384
rect 844 1376 852 1384
rect 940 1376 948 1384
rect 1164 1376 1172 1384
rect 1212 1376 1220 1384
rect 1292 1376 1300 1384
rect 1980 1376 1988 1384
rect 236 1356 244 1364
rect 556 1356 564 1364
rect 716 1356 724 1364
rect 780 1356 788 1364
rect 860 1356 868 1364
rect 1372 1356 1380 1364
rect 1548 1356 1556 1364
rect 1852 1356 1860 1364
rect 2188 1356 2196 1364
rect 268 1336 276 1344
rect 412 1336 420 1344
rect 828 1336 836 1344
rect 876 1336 884 1344
rect 972 1336 980 1344
rect 1052 1336 1060 1344
rect 1276 1336 1284 1344
rect 1516 1336 1524 1344
rect 1900 1336 1908 1344
rect 1916 1336 1924 1344
rect 2012 1336 2020 1344
rect 2156 1336 2164 1344
rect 2350 1336 2358 1344
rect 44 1316 52 1324
rect 268 1316 276 1324
rect 380 1316 388 1324
rect 524 1316 532 1324
rect 604 1316 612 1324
rect 636 1316 644 1324
rect 652 1316 660 1324
rect 812 1316 820 1324
rect 828 1316 836 1324
rect 988 1316 996 1324
rect 1196 1316 1204 1324
rect 1324 1316 1332 1324
rect 1420 1316 1428 1324
rect 1788 1316 1796 1324
rect 1820 1316 1828 1324
rect 2092 1316 2100 1324
rect 364 1296 372 1304
rect 588 1296 596 1304
rect 1244 1296 1252 1304
rect 1292 1296 1300 1304
rect 1452 1300 1460 1308
rect 1708 1296 1716 1304
rect 1852 1296 1860 1304
rect 2060 1296 2068 1304
rect 12 1276 20 1284
rect 60 1276 68 1284
rect 668 1276 676 1284
rect 652 1256 660 1264
rect 1020 1256 1028 1264
rect 364 1236 372 1244
rect 572 1236 580 1244
rect 1452 1236 1460 1244
rect 1884 1236 1892 1244
rect 2060 1236 2068 1244
rect 686 1206 694 1214
rect 700 1206 708 1214
rect 714 1206 722 1214
rect 364 1176 372 1184
rect 812 1176 820 1184
rect 1244 1176 1252 1184
rect 1292 1176 1300 1184
rect 1356 1176 1364 1184
rect 1900 1176 1908 1184
rect 2252 1176 2260 1184
rect 2396 1176 2404 1184
rect 76 1136 84 1144
rect 828 1136 836 1144
rect 908 1136 916 1144
rect 940 1136 948 1144
rect 1164 1136 1172 1144
rect 1180 1136 1188 1144
rect 1276 1136 1284 1144
rect 1644 1136 1652 1144
rect 1820 1136 1828 1144
rect 2300 1136 2308 1144
rect 364 1116 372 1124
rect 524 1116 532 1124
rect 796 1116 804 1124
rect 972 1116 980 1124
rect 1052 1116 1060 1124
rect 1148 1116 1156 1124
rect 1308 1116 1316 1124
rect 1356 1116 1364 1124
rect 1756 1116 1764 1124
rect 1900 1116 1908 1124
rect 268 1096 276 1104
rect 364 1096 372 1104
rect 604 1096 612 1104
rect 748 1096 756 1104
rect 812 1096 820 1104
rect 892 1096 900 1104
rect 956 1096 964 1104
rect 1020 1096 1028 1104
rect 1132 1096 1140 1104
rect 1164 1096 1172 1104
rect 1244 1096 1252 1104
rect 1292 1096 1300 1104
rect 1372 1096 1380 1104
rect 1564 1096 1572 1104
rect 1900 1096 1908 1104
rect 2108 1096 2116 1104
rect 2268 1096 2276 1104
rect 2316 1096 2324 1104
rect 2364 1096 2372 1104
rect 12 1076 20 1084
rect 268 1076 276 1084
rect 412 1076 420 1084
rect 508 1076 516 1084
rect 540 1076 548 1084
rect 556 1076 564 1084
rect 748 1076 756 1084
rect 1036 1076 1044 1084
rect 1084 1076 1092 1084
rect 1452 1076 1460 1084
rect 1660 1076 1668 1084
rect 1772 1076 1780 1084
rect 1852 1076 1860 1084
rect 1996 1076 2004 1084
rect 2348 1076 2356 1084
rect 236 1056 244 1064
rect 572 1056 580 1064
rect 620 1056 628 1064
rect 748 1056 756 1064
rect 860 1056 868 1064
rect 892 1056 900 1064
rect 1100 1056 1108 1064
rect 1212 1056 1220 1064
rect 1484 1056 1492 1064
rect 2028 1056 2036 1064
rect 444 1036 452 1044
rect 588 1036 596 1044
rect 748 1036 756 1044
rect 956 1036 964 1044
rect 988 1036 996 1044
rect 1052 1036 1060 1044
rect 1164 1036 1172 1044
rect 2188 1036 2196 1044
rect 1694 1006 1702 1014
rect 1708 1006 1716 1014
rect 1722 1006 1730 1014
rect 172 976 180 984
rect 396 976 404 984
rect 524 976 532 984
rect 732 976 740 984
rect 780 976 788 984
rect 1004 976 1012 984
rect 1212 976 1220 984
rect 1292 976 1300 984
rect 1436 976 1444 984
rect 1532 976 1540 984
rect 1964 976 1972 984
rect 492 956 500 964
rect 572 956 580 964
rect 588 956 596 964
rect 748 956 756 964
rect 892 956 900 964
rect 908 956 916 964
rect 1020 956 1028 964
rect 1084 956 1092 964
rect 1132 956 1140 964
rect 1340 956 1348 964
rect 1452 956 1460 964
rect 1580 956 1588 964
rect 1788 956 1796 964
rect 1900 956 1908 964
rect 2140 956 2148 964
rect 2316 956 2324 964
rect 12 936 20 944
rect 60 936 68 944
rect 332 936 340 944
rect 348 936 356 944
rect 444 936 452 944
rect 460 936 468 944
rect 1052 936 1060 944
rect 1100 936 1108 944
rect 1132 936 1140 944
rect 1196 936 1204 944
rect 1244 936 1252 944
rect 1260 936 1268 944
rect 1292 936 1300 944
rect 1484 936 1492 944
rect 1724 936 1732 944
rect 1916 936 1924 944
rect 2108 936 2116 944
rect 44 916 52 924
rect 460 916 468 924
rect 556 916 564 924
rect 620 916 628 924
rect 780 916 788 924
rect 844 916 852 924
rect 988 916 996 924
rect 1052 916 1060 924
rect 1100 916 1108 924
rect 1228 916 1236 924
rect 1420 916 1428 924
rect 1580 916 1588 924
rect 1644 916 1652 924
rect 1740 916 1748 924
rect 1788 916 1796 924
rect 1836 916 1844 924
rect 1868 916 1876 924
rect 1932 916 1940 924
rect 2028 916 2036 924
rect 2316 916 2324 924
rect 604 896 612 904
rect 764 896 772 904
rect 828 896 836 904
rect 1116 896 1124 904
rect 1180 896 1188 904
rect 1532 896 1540 904
rect 1596 896 1604 904
rect 1660 896 1668 904
rect 2044 900 2052 908
rect 636 876 644 884
rect 796 876 804 884
rect 860 876 868 884
rect 1196 876 1204 884
rect 1564 876 1572 884
rect 1596 876 1604 884
rect 1628 876 1636 884
rect 780 856 788 864
rect 1724 876 1732 884
rect 2396 876 2404 884
rect 2044 854 2052 862
rect 220 836 228 844
rect 876 836 884 844
rect 2300 836 2308 844
rect 686 806 694 814
rect 700 806 708 814
rect 714 806 722 814
rect 364 776 372 784
rect 716 776 724 784
rect 1132 776 1140 784
rect 1292 776 1300 784
rect 1628 776 1636 784
rect 876 758 884 766
rect 1548 758 1556 766
rect 2044 758 2052 766
rect 12 736 20 744
rect 1772 736 1780 744
rect 2316 736 2324 744
rect 364 716 372 724
rect 716 716 724 724
rect 876 712 884 720
rect 1548 712 1556 720
rect 1676 716 1684 724
rect 1804 716 1812 724
rect 2044 712 2052 720
rect 364 696 372 704
rect 508 696 516 704
rect 716 696 724 704
rect 1052 696 1060 704
rect 1276 696 1284 704
rect 1564 696 1572 704
rect 1660 696 1668 704
rect 1788 696 1796 704
rect 1852 696 1860 704
rect 1964 696 1972 704
rect 2028 696 2036 704
rect 2302 696 2310 704
rect 2332 696 2340 704
rect 268 676 276 684
rect 620 676 628 684
rect 940 676 948 684
rect 1484 676 1492 684
rect 1772 676 1780 684
rect 1884 676 1892 684
rect 1964 676 1972 684
rect 2108 676 2116 684
rect 2396 676 2404 684
rect 236 656 244 664
rect 588 656 596 664
rect 972 656 980 664
rect 1452 656 1460 664
rect 1644 656 1652 664
rect 1692 656 1700 664
rect 1820 656 1828 664
rect 1852 656 1860 664
rect 1868 656 1876 664
rect 1932 656 1940 664
rect 2140 656 2148 664
rect 76 636 84 644
rect 428 636 436 644
rect 1132 636 1140 644
rect 1916 636 1924 644
rect 1694 606 1702 614
rect 1708 606 1716 614
rect 1722 606 1730 614
rect 316 576 324 584
rect 620 576 628 584
rect 812 576 820 584
rect 956 576 964 584
rect 1116 576 1124 584
rect 1148 576 1156 584
rect 1212 576 1220 584
rect 1868 576 1876 584
rect 108 556 116 564
rect 124 556 132 564
rect 188 556 196 564
rect 204 556 212 564
rect 60 536 68 544
rect 140 536 148 544
rect 236 536 244 544
rect 268 536 276 544
rect 364 536 372 544
rect 380 536 388 544
rect 460 536 468 544
rect 492 536 500 544
rect 588 536 596 544
rect 652 556 660 564
rect 972 556 980 564
rect 1004 556 1012 564
rect 1036 556 1044 564
rect 1132 556 1140 564
rect 1436 556 1444 564
rect 1884 556 1892 564
rect 1980 556 1988 564
rect 2172 556 2180 564
rect 716 536 724 544
rect 844 532 852 540
rect 860 536 868 544
rect 876 536 884 544
rect 908 536 916 544
rect 1100 536 1108 544
rect 1180 532 1188 540
rect 1244 536 1252 544
rect 1468 536 1476 544
rect 1612 536 1620 544
rect 1740 536 1748 544
rect 1788 536 1796 544
rect 1948 536 1956 544
rect 1996 536 2004 544
rect 2140 536 2148 544
rect 220 516 228 524
rect 252 516 260 524
rect 364 516 372 524
rect 604 516 612 524
rect 748 516 756 524
rect 796 516 804 524
rect 924 516 932 524
rect 1004 516 1012 524
rect 1052 516 1060 524
rect 1068 516 1076 524
rect 1564 516 1572 524
rect 1932 516 1940 524
rect 2044 516 2052 524
rect 76 496 84 504
rect 92 496 100 504
rect 428 496 436 504
rect 556 496 564 504
rect 908 496 916 504
rect 972 496 980 504
rect 1212 496 1220 504
rect 1532 500 1540 508
rect 1836 496 1844 504
rect 1900 496 1908 504
rect 1932 496 1940 504
rect 1964 496 1972 504
rect 2076 500 2084 508
rect 12 476 20 484
rect 540 476 548 484
rect 1244 476 1252 484
rect 1532 454 1540 462
rect 2076 454 2084 462
rect 572 436 580 444
rect 2332 436 2340 444
rect 686 406 694 414
rect 700 406 708 414
rect 714 406 722 414
rect 28 376 36 384
rect 316 376 324 384
rect 444 376 452 384
rect 972 376 980 384
rect 1996 376 2004 384
rect 2108 376 2116 384
rect 1548 358 1556 366
rect 2124 336 2132 344
rect 316 316 324 324
rect 444 316 452 324
rect 956 316 964 324
rect 1020 316 1028 324
rect 1548 312 1556 320
rect 2012 316 2020 324
rect 316 296 324 304
rect 396 296 404 304
rect 476 296 484 304
rect 652 296 660 304
rect 748 296 756 304
rect 220 276 228 284
rect 540 276 548 284
rect 812 276 820 284
rect 924 296 932 304
rect 1100 296 1108 304
rect 1116 296 1124 304
rect 1180 296 1188 304
rect 1260 296 1268 304
rect 1564 296 1572 304
rect 1580 296 1588 304
rect 1852 296 1860 304
rect 2044 296 2052 304
rect 2108 296 2116 304
rect 2156 296 2164 304
rect 2220 296 2228 304
rect 2284 296 2292 304
rect 2332 296 2340 304
rect 924 276 932 284
rect 1068 276 1076 284
rect 1132 280 1140 288
rect 188 256 196 264
rect 572 256 580 264
rect 1068 256 1076 264
rect 1212 256 1220 264
rect 1290 276 1298 284
rect 1484 276 1492 284
rect 1676 276 1684 284
rect 1868 276 1876 284
rect 1980 276 1988 284
rect 2172 276 2180 284
rect 2236 276 2244 284
rect 2252 276 2260 284
rect 2316 276 2324 284
rect 1276 256 1284 264
rect 1452 256 1460 264
rect 1788 256 1796 264
rect 2060 256 2068 264
rect 2204 256 2212 264
rect 2268 256 2276 264
rect 364 236 372 244
rect 1164 236 1172 244
rect 1820 236 1828 244
rect 1900 236 1908 244
rect 2188 236 2196 244
rect 2364 236 2372 244
rect 1694 206 1702 214
rect 1708 206 1716 214
rect 1722 206 1730 214
rect 28 176 36 184
rect 892 176 900 184
rect 1036 176 1044 184
rect 1324 176 1332 184
rect 1484 176 1492 184
rect 1580 176 1588 184
rect 1980 176 1988 184
rect 2332 176 2340 184
rect 188 156 196 164
rect 732 156 740 164
rect 1020 156 1028 164
rect 1052 156 1060 164
rect 1100 156 1108 164
rect 1820 156 1828 164
rect 2172 156 2180 164
rect 220 136 228 144
rect 412 136 420 144
rect 508 136 516 144
rect 700 136 708 144
rect 1132 136 1140 144
rect 1260 136 1268 144
rect 1356 136 1364 144
rect 1532 136 1540 144
rect 1788 136 1796 144
rect 2140 136 2148 144
rect 316 116 324 124
rect 364 116 372 124
rect 412 116 420 124
rect 620 116 628 124
rect 924 116 932 124
rect 972 116 980 124
rect 1052 116 1060 124
rect 1148 116 1156 124
rect 1196 116 1204 124
rect 1212 116 1220 124
rect 1420 116 1428 124
rect 1692 116 1700 124
rect 1900 116 1908 124
rect 2044 116 2052 124
rect 284 100 292 108
rect 636 100 644 108
rect 1724 100 1732 108
rect 2076 100 2084 108
rect 1724 54 1732 62
rect 2076 54 2084 62
rect 284 36 292 44
rect 396 36 404 44
rect 636 36 644 44
rect 956 36 964 44
rect 1004 36 1012 44
rect 1164 36 1172 44
rect 1244 36 1252 44
rect 1404 36 1412 44
rect 1452 36 1460 44
rect 686 6 694 14
rect 700 6 708 14
rect 714 6 722 14
<< metal2 >>
rect 381 2037 403 2043
rect 429 2037 451 2043
rect 397 1984 403 2037
rect 445 1984 451 2037
rect 680 2006 686 2014
rect 694 2006 700 2014
rect 708 2006 714 2014
rect 722 2006 728 2014
rect 781 2004 787 2043
rect 861 2037 883 2043
rect 1293 2037 1315 2043
rect 1341 2037 1363 2043
rect 1485 2037 1507 2043
rect 1853 2037 1875 2043
rect 1997 2037 2019 2043
rect 861 1984 867 2037
rect 1309 1984 1315 2037
rect 1357 1984 1363 2037
rect 317 1924 323 1976
rect 493 1924 499 1976
rect 372 1897 387 1903
rect 317 1884 323 1896
rect 29 1784 35 1836
rect 77 1784 83 1876
rect 13 1777 28 1783
rect 13 1744 19 1777
rect 189 1764 195 1856
rect 157 1644 163 1696
rect 189 1464 195 1756
rect 253 1724 259 1736
rect 365 1724 371 1876
rect 381 1784 387 1897
rect 413 1804 419 1896
rect 493 1884 499 1896
rect 589 1844 595 1876
rect 445 1784 451 1796
rect 589 1744 595 1776
rect 317 1524 323 1576
rect 365 1504 371 1716
rect 397 1524 403 1576
rect 388 1497 396 1503
rect 29 1323 35 1436
rect 189 1424 195 1456
rect 221 1404 227 1476
rect 237 1364 243 1416
rect 29 1317 44 1323
rect 13 1284 19 1296
rect 13 1084 19 1096
rect 61 984 67 1276
rect 77 1124 83 1136
rect 237 1064 243 1356
rect 381 1324 387 1496
rect 493 1484 499 1516
rect 525 1424 531 1456
rect 621 1424 627 1856
rect 653 1744 659 1756
rect 701 1744 707 1876
rect 717 1744 723 1796
rect 781 1784 787 1936
rect 1469 1924 1475 1976
rect 957 1917 972 1923
rect 877 1897 892 1903
rect 653 1724 659 1736
rect 445 1384 451 1396
rect 269 1104 275 1316
rect 365 1244 371 1296
rect 237 1024 243 1056
rect 269 1044 275 1076
rect 173 984 179 1016
rect 13 904 19 936
rect 45 924 51 976
rect 333 964 339 1176
rect 365 1124 371 1176
rect 397 984 403 1336
rect 557 1284 563 1356
rect 589 1304 595 1336
rect 637 1324 643 1496
rect 653 1344 659 1716
rect 749 1704 755 1776
rect 813 1744 819 1856
rect 680 1606 686 1614
rect 694 1606 700 1614
rect 708 1606 714 1614
rect 722 1606 728 1614
rect 765 1584 771 1696
rect 605 1304 611 1316
rect 653 1304 659 1316
rect 669 1284 675 1536
rect 717 1464 723 1576
rect 829 1544 835 1636
rect 877 1584 883 1897
rect 909 1804 915 1876
rect 925 1784 931 1896
rect 957 1784 963 1917
rect 1005 1884 1011 1896
rect 973 1763 979 1836
rect 1085 1784 1091 1836
rect 1101 1824 1107 1896
rect 1165 1884 1171 1896
rect 1197 1884 1203 1916
rect 1261 1904 1267 1916
rect 1389 1904 1395 1916
rect 1213 1844 1219 1876
rect 1261 1864 1267 1896
rect 1101 1764 1107 1816
rect 1293 1764 1299 1856
rect 1325 1824 1331 1896
rect 1469 1884 1475 1896
rect 1373 1864 1379 1876
rect 1405 1824 1411 1876
rect 957 1757 979 1763
rect 925 1704 931 1716
rect 916 1697 924 1703
rect 717 1364 723 1456
rect 717 1304 723 1356
rect 653 1264 659 1276
rect 669 1244 675 1276
rect 413 1084 419 1116
rect 509 1044 515 1076
rect 525 984 531 1096
rect 557 984 563 1076
rect 573 1064 579 1236
rect 680 1206 686 1214
rect 694 1206 700 1214
rect 708 1206 714 1214
rect 722 1206 728 1214
rect 61 944 67 956
rect 333 944 339 956
rect 445 944 451 976
rect 589 964 595 1036
rect 461 884 467 916
rect 605 904 611 976
rect 621 924 627 1056
rect 637 884 643 1016
rect 669 924 675 1156
rect 749 1104 755 1376
rect 781 1364 787 1476
rect 909 1444 915 1476
rect 845 1384 851 1436
rect 941 1384 947 1476
rect 957 1384 963 1757
rect 1069 1724 1075 1736
rect 861 1364 867 1376
rect 973 1344 979 1496
rect 989 1324 995 1496
rect 1101 1464 1107 1676
rect 1213 1504 1219 1716
rect 1293 1684 1299 1756
rect 1437 1724 1443 1876
rect 1501 1784 1507 2037
rect 1869 1984 1875 2037
rect 2013 1984 2019 2037
rect 2061 1924 2067 1976
rect 1565 1884 1571 1916
rect 1933 1904 1939 1916
rect 1933 1884 1939 1896
rect 1853 1844 1859 1856
rect 1517 1784 1523 1816
rect 1688 1806 1694 1814
rect 1702 1806 1708 1814
rect 1716 1806 1722 1814
rect 1730 1806 1736 1814
rect 1581 1764 1587 1776
rect 1757 1764 1763 1836
rect 1437 1704 1443 1716
rect 1389 1662 1395 1700
rect 1357 1584 1363 1616
rect 1229 1524 1235 1576
rect 1437 1504 1443 1696
rect 1469 1624 1475 1716
rect 1597 1704 1603 1756
rect 1821 1744 1827 1796
rect 1853 1764 1859 1836
rect 1933 1784 1939 1836
rect 1549 1524 1555 1636
rect 1677 1584 1683 1736
rect 1725 1704 1731 1716
rect 1933 1703 1939 1716
rect 1949 1703 1955 1876
rect 1965 1784 1971 1876
rect 2013 1784 2019 1896
rect 2061 1884 2067 1896
rect 2157 1823 2163 1876
rect 2189 1844 2195 1856
rect 2157 1817 2179 1823
rect 2077 1784 2083 1796
rect 2173 1784 2179 1817
rect 1757 1662 1763 1700
rect 1933 1697 1955 1703
rect 1645 1524 1651 1576
rect 1949 1504 1955 1697
rect 2157 1524 2163 1576
rect 1229 1484 1235 1496
rect 1853 1484 1859 1496
rect 1101 1424 1107 1456
rect 1165 1384 1171 1416
rect 1213 1384 1219 1456
rect 1293 1384 1299 1476
rect 1517 1444 1523 1456
rect 1741 1444 1747 1476
rect 1364 1437 1379 1443
rect 1373 1364 1379 1437
rect 1549 1364 1555 1436
rect 1688 1406 1694 1414
rect 1702 1406 1708 1414
rect 1716 1406 1722 1414
rect 1730 1406 1736 1414
rect 733 984 739 1036
rect 749 984 755 1036
rect 765 923 771 1036
rect 781 984 787 1316
rect 813 1184 819 1316
rect 941 1144 947 1236
rect 989 1164 995 1316
rect 1053 1184 1059 1336
rect 1325 1324 1331 1336
rect 797 1044 803 1116
rect 813 1104 819 1116
rect 829 1024 835 1136
rect 941 1124 947 1136
rect 973 1124 979 1136
rect 1021 1104 1027 1116
rect 1037 1084 1043 1156
rect 893 1064 899 1076
rect 749 917 771 923
rect 669 844 675 916
rect 221 783 227 836
rect 680 806 686 814
rect 694 806 700 814
rect 708 806 714 814
rect 722 806 728 814
rect 221 777 243 783
rect 13 704 19 736
rect 237 664 243 777
rect 365 724 371 776
rect 717 724 723 776
rect 13 484 19 496
rect 29 384 35 556
rect 61 544 67 556
rect 77 543 83 636
rect 269 624 275 676
rect 189 564 195 576
rect 253 564 259 596
rect 317 584 323 616
rect 77 537 92 543
rect 93 504 99 536
rect 237 524 243 536
rect 253 524 259 556
rect 301 550 307 576
rect 381 524 387 536
rect 429 524 435 636
rect 221 284 227 516
rect 365 504 371 516
rect 317 324 323 376
rect 397 304 403 516
rect 429 504 435 516
rect 445 324 451 376
rect 189 164 195 256
rect 221 124 227 136
rect 317 124 323 296
rect 372 237 387 243
rect 365 124 371 176
rect 285 44 291 100
rect 381 -23 387 237
rect 461 184 467 536
rect 477 304 483 696
rect 621 584 627 676
rect 589 544 595 556
rect 717 544 723 696
rect 749 544 755 917
rect 765 904 771 917
rect 797 884 803 996
rect 845 924 851 996
rect 813 903 819 916
rect 813 897 828 903
rect 781 864 787 876
rect 557 504 563 536
rect 589 524 595 536
rect 749 524 755 536
rect 797 524 803 836
rect 813 584 819 897
rect 861 884 867 976
rect 909 964 915 1036
rect 957 924 963 1036
rect 989 1004 995 1036
rect 1005 884 1011 976
rect 1053 944 1059 1036
rect 1053 924 1059 936
rect 877 720 883 758
rect 1069 703 1075 1256
rect 1085 1084 1091 1156
rect 1133 1104 1139 1316
rect 1149 1124 1155 1136
rect 1085 964 1091 996
rect 1060 697 1075 703
rect 941 644 947 676
rect 1085 624 1091 956
rect 1101 944 1107 1016
rect 1133 1004 1139 1096
rect 1165 1063 1171 1096
rect 1181 1084 1187 1136
rect 1165 1057 1187 1063
rect 1165 964 1171 1036
rect 1181 1004 1187 1057
rect 1197 944 1203 1296
rect 1245 1184 1251 1296
rect 1293 1184 1299 1276
rect 1245 1164 1251 1176
rect 1325 1124 1331 1316
rect 1421 1264 1427 1316
rect 1293 1104 1299 1116
rect 1213 984 1219 1056
rect 1245 944 1251 1016
rect 1293 984 1299 1056
rect 1309 1024 1315 1116
rect 1325 1044 1331 1116
rect 1341 964 1347 1136
rect 1357 1124 1363 1176
rect 1373 1104 1379 1256
rect 1453 1244 1459 1300
rect 1549 1224 1555 1356
rect 1773 1344 1779 1436
rect 1789 1324 1795 1436
rect 1853 1364 1859 1476
rect 2029 1444 2035 1456
rect 2189 1444 2195 1836
rect 2381 1784 2387 1856
rect 2205 1764 2211 1776
rect 2381 1764 2387 1776
rect 2205 1504 2211 1736
rect 2237 1724 2243 1736
rect 2253 1584 2259 1736
rect 2333 1724 2339 1756
rect 2269 1697 2284 1703
rect 2253 1464 2259 1496
rect 2269 1463 2275 1697
rect 2285 1464 2291 1576
rect 2349 1504 2355 1576
rect 2333 1484 2339 1496
rect 2260 1457 2275 1463
rect 1789 1284 1795 1316
rect 1853 1304 1859 1356
rect 2157 1344 2163 1376
rect 2189 1364 2195 1436
rect 1917 1324 1923 1336
rect 2061 1244 2067 1296
rect 1453 1064 1459 1076
rect 1485 1064 1491 1216
rect 1565 1064 1571 1096
rect 1485 1023 1491 1056
rect 1469 1017 1491 1023
rect 1229 924 1235 936
rect 1197 784 1203 876
rect 1245 784 1251 936
rect 1261 904 1267 936
rect 1293 864 1299 936
rect 1437 924 1443 976
rect 1453 944 1459 956
rect 1421 844 1427 916
rect 1469 903 1475 1017
rect 1485 944 1491 976
rect 1533 904 1539 936
rect 1645 924 1651 996
rect 1661 944 1667 1076
rect 1688 1006 1694 1014
rect 1702 1006 1708 1014
rect 1716 1006 1722 1014
rect 1730 1006 1736 1014
rect 1725 944 1731 976
rect 1453 897 1475 903
rect 1277 684 1283 696
rect 957 584 963 616
rect 1117 584 1123 676
rect 1453 664 1459 897
rect 1533 844 1539 896
rect 1565 884 1571 896
rect 1581 864 1587 916
rect 1629 884 1635 916
rect 1661 904 1667 936
rect 1741 924 1747 956
rect 1629 784 1635 836
rect 1549 720 1555 758
rect 1645 744 1651 896
rect 1133 564 1139 636
rect 1149 584 1155 636
rect 1213 584 1219 664
rect 1453 623 1459 656
rect 1437 617 1459 623
rect 1437 564 1443 617
rect 845 540 851 556
rect 605 484 611 516
rect 541 284 547 296
rect 573 284 579 436
rect 680 406 686 414
rect 694 406 700 414
rect 708 406 714 414
rect 722 406 728 414
rect 653 204 659 296
rect 413 144 419 176
rect 621 124 627 196
rect 733 164 739 256
rect 797 204 803 516
rect 861 504 867 536
rect 909 504 915 536
rect 925 304 931 516
rect 973 504 979 556
rect 1053 504 1059 516
rect 973 384 979 496
rect 813 164 819 276
rect 925 184 931 276
rect 957 184 963 316
rect 893 144 899 176
rect 1021 164 1027 316
rect 1037 184 1043 256
rect 1053 164 1059 496
rect 1101 304 1107 516
rect 701 124 707 136
rect 925 124 931 156
rect 1101 144 1107 156
rect 1133 144 1139 176
rect 1165 144 1171 236
rect 973 124 979 136
rect 1165 123 1171 136
rect 1197 124 1203 556
rect 1245 544 1251 556
rect 1213 264 1219 276
rect 1213 124 1219 256
rect 1245 184 1251 476
rect 1261 144 1267 296
rect 1325 184 1331 536
rect 1437 443 1443 556
rect 1565 524 1571 696
rect 1645 664 1651 736
rect 1661 704 1667 876
rect 1757 864 1763 1116
rect 1885 1104 1891 1236
rect 2093 1223 2099 1316
rect 2093 1217 2115 1223
rect 1901 1124 1907 1176
rect 2109 1104 2115 1217
rect 2269 1104 2275 1136
rect 1805 943 1811 956
rect 1789 937 1811 943
rect 1789 924 1795 937
rect 1757 743 1763 856
rect 1853 844 1859 1076
rect 1901 1064 1907 1096
rect 1901 964 1907 1036
rect 1997 1024 2003 1076
rect 1965 984 1971 1016
rect 2109 1004 2115 1096
rect 1901 944 1907 956
rect 1917 884 1923 936
rect 2029 924 2035 996
rect 2141 964 2147 1056
rect 2317 964 2323 1096
rect 2109 944 2115 956
rect 1805 744 1811 836
rect 1757 737 1772 743
rect 1805 724 1811 736
rect 1853 704 1859 816
rect 1965 704 1971 716
rect 2029 704 2035 916
rect 2045 862 2051 900
rect 2045 720 2051 758
rect 1789 664 1795 696
rect 1853 683 1859 696
rect 1853 677 1875 683
rect 1821 664 1827 676
rect 1869 664 1875 677
rect 2141 664 2147 956
rect 2317 744 2323 916
rect 2333 704 2339 1336
rect 2381 1103 2387 1756
rect 2397 1184 2403 1216
rect 2372 1097 2387 1103
rect 2349 1084 2355 1096
rect 2397 884 2403 896
rect 2397 684 2403 696
rect 1688 606 1694 614
rect 1702 606 1708 614
rect 1716 606 1722 614
rect 1730 606 1736 614
rect 1789 544 1795 656
rect 1533 462 1539 500
rect 1437 437 1459 443
rect 1453 264 1459 437
rect 1549 320 1555 358
rect 1565 304 1571 516
rect 1485 184 1491 196
rect 1581 184 1587 296
rect 1677 284 1683 536
rect 1837 303 1843 496
rect 1853 323 1859 656
rect 1869 584 1875 636
rect 1885 464 1891 556
rect 1917 523 1923 636
rect 2141 624 2147 656
rect 2173 564 2179 616
rect 2141 544 2147 556
rect 2173 544 2179 556
rect 2004 537 2019 543
rect 1917 517 1932 523
rect 1949 464 1955 536
rect 1997 384 2003 456
rect 2013 424 2019 537
rect 2029 517 2044 523
rect 1869 323 1875 336
rect 1853 317 1875 323
rect 1837 297 1852 303
rect 1853 284 1859 296
rect 1869 284 1875 317
rect 1981 264 1987 276
rect 1688 206 1694 214
rect 1702 206 1708 214
rect 1716 206 1722 214
rect 1730 206 1736 214
rect 1821 184 1827 236
rect 1357 144 1363 176
rect 1156 117 1171 123
rect 637 44 643 100
rect 1533 44 1539 136
rect 1581 124 1587 176
rect 1901 144 1907 236
rect 1981 184 1987 256
rect 2029 124 2035 517
rect 2077 462 2083 500
rect 2061 284 2067 436
rect 2109 384 2115 416
rect 2173 284 2179 336
rect 2221 304 2227 336
rect 2061 264 2067 276
rect 2205 264 2211 276
rect 2237 264 2243 276
rect 2269 264 2275 316
rect 2333 304 2339 316
rect 2285 264 2291 296
rect 2317 284 2323 296
rect 2141 144 2147 196
rect 2173 164 2179 216
rect 2189 204 2195 236
rect 2333 184 2339 296
rect 1725 62 1731 100
rect 2077 62 2083 100
rect 397 -17 403 36
rect 957 24 963 36
rect 680 6 686 14
rect 694 6 700 14
rect 708 6 714 14
rect 722 6 728 14
rect 397 -23 419 -17
rect 925 -23 931 16
rect 1005 -17 1011 36
rect 989 -23 1011 -17
rect 1165 -17 1171 36
rect 1245 -17 1251 36
rect 1405 -17 1411 36
rect 1453 -17 1459 36
rect 1165 -23 1187 -17
rect 1229 -23 1251 -17
rect 1389 -23 1411 -17
rect 1437 -23 1459 -17
rect 1501 -23 1507 36
rect 1837 -23 1843 16
rect 2365 -17 2371 236
rect 2349 -23 2371 -17
<< m3contact >>
rect 686 2006 694 2014
rect 700 2006 708 2014
rect 714 2006 722 2014
rect 780 1996 788 2004
rect 780 1936 788 1944
rect 1084 1936 1092 1944
rect 76 1876 84 1884
rect 220 1876 228 1884
rect 316 1876 324 1884
rect 364 1876 372 1884
rect 28 1776 36 1784
rect 188 1756 196 1764
rect 284 1756 292 1764
rect 108 1736 116 1744
rect 492 1876 500 1884
rect 700 1876 708 1884
rect 588 1836 596 1844
rect 412 1796 420 1804
rect 444 1796 452 1804
rect 380 1776 388 1784
rect 588 1776 596 1784
rect 252 1716 260 1724
rect 460 1716 468 1724
rect 492 1516 500 1524
rect 316 1496 324 1504
rect 364 1496 372 1504
rect 380 1496 388 1504
rect 188 1416 196 1424
rect 236 1416 244 1424
rect 220 1396 228 1404
rect 44 1316 52 1324
rect 12 1296 20 1304
rect 12 1096 20 1104
rect 76 1116 84 1124
rect 268 1336 276 1344
rect 716 1796 724 1804
rect 812 1856 820 1864
rect 748 1776 756 1784
rect 652 1736 660 1744
rect 652 1716 660 1724
rect 636 1496 644 1504
rect 524 1416 532 1424
rect 620 1416 628 1424
rect 444 1396 452 1404
rect 396 1336 404 1344
rect 412 1336 420 1344
rect 332 1176 340 1184
rect 268 1036 276 1044
rect 172 1016 180 1024
rect 236 1016 244 1024
rect 44 976 52 984
rect 60 976 68 984
rect 364 1096 372 1104
rect 524 1316 532 1324
rect 588 1336 596 1344
rect 764 1756 772 1764
rect 796 1756 804 1764
rect 812 1736 820 1744
rect 860 1736 868 1744
rect 764 1716 772 1724
rect 764 1696 772 1704
rect 686 1606 694 1614
rect 700 1606 708 1614
rect 714 1606 722 1614
rect 716 1576 724 1584
rect 668 1536 676 1544
rect 652 1336 660 1344
rect 604 1296 612 1304
rect 652 1296 660 1304
rect 908 1796 916 1804
rect 1020 1916 1028 1924
rect 1228 1916 1236 1924
rect 1388 1916 1396 1924
rect 972 1896 980 1904
rect 1004 1896 1012 1904
rect 1164 1896 1172 1904
rect 1020 1836 1028 1844
rect 1084 1836 1092 1844
rect 924 1776 932 1784
rect 1420 1896 1428 1904
rect 1196 1876 1204 1884
rect 1148 1856 1156 1864
rect 1260 1856 1268 1864
rect 1292 1856 1300 1864
rect 1212 1836 1220 1844
rect 1100 1816 1108 1824
rect 1372 1876 1380 1884
rect 1436 1876 1444 1884
rect 1468 1876 1476 1884
rect 1324 1816 1332 1824
rect 1404 1816 1412 1824
rect 892 1736 900 1744
rect 924 1696 932 1704
rect 876 1576 884 1584
rect 828 1536 836 1544
rect 844 1516 852 1524
rect 796 1496 804 1504
rect 940 1496 946 1504
rect 946 1496 948 1504
rect 780 1476 788 1484
rect 812 1476 820 1484
rect 940 1476 948 1484
rect 748 1376 756 1384
rect 716 1296 724 1304
rect 556 1276 564 1284
rect 652 1276 660 1284
rect 668 1236 676 1244
rect 412 1116 420 1124
rect 524 1116 532 1124
rect 524 1096 532 1104
rect 444 1036 452 1044
rect 508 1036 516 1044
rect 540 1076 548 1084
rect 686 1206 694 1214
rect 700 1206 708 1214
rect 714 1206 722 1214
rect 668 1156 676 1164
rect 604 1096 612 1104
rect 572 1056 580 1064
rect 444 976 452 984
rect 556 976 564 984
rect 60 956 68 964
rect 332 956 340 964
rect 604 976 612 984
rect 492 956 500 964
rect 572 956 580 964
rect 348 936 356 944
rect 460 936 468 944
rect 556 916 564 924
rect 12 896 20 904
rect 636 1016 644 1024
rect 844 1436 852 1444
rect 908 1436 916 1444
rect 972 1736 980 1744
rect 1068 1736 1076 1744
rect 1116 1696 1124 1704
rect 1100 1676 1108 1684
rect 972 1496 980 1504
rect 988 1496 996 1504
rect 860 1376 868 1384
rect 956 1376 964 1384
rect 828 1336 836 1344
rect 876 1336 884 1344
rect 1324 1736 1332 1744
rect 1564 1916 1572 1924
rect 1884 1916 1892 1924
rect 1884 1896 1892 1904
rect 1932 1896 1940 1904
rect 1980 1896 1988 1904
rect 2012 1896 2020 1904
rect 1948 1876 1956 1884
rect 1596 1856 1604 1864
rect 1852 1856 1860 1864
rect 1852 1836 1860 1844
rect 1516 1816 1524 1824
rect 1694 1806 1702 1814
rect 1708 1806 1716 1814
rect 1722 1806 1730 1814
rect 1580 1776 1588 1784
rect 1820 1796 1828 1804
rect 1532 1756 1540 1764
rect 1596 1756 1604 1764
rect 1756 1756 1764 1764
rect 1548 1716 1556 1724
rect 1580 1716 1588 1724
rect 1292 1676 1300 1684
rect 1436 1696 1444 1704
rect 1356 1616 1364 1624
rect 1932 1776 1940 1784
rect 1468 1616 1476 1624
rect 1724 1696 1732 1704
rect 2060 1876 2068 1884
rect 2188 1836 2196 1844
rect 2076 1796 2084 1804
rect 1964 1776 1972 1784
rect 2156 1756 2164 1764
rect 1676 1576 1684 1584
rect 1868 1576 1876 1584
rect 1548 1516 1556 1524
rect 1324 1496 1332 1504
rect 1852 1496 1860 1504
rect 1132 1476 1140 1484
rect 1228 1476 1236 1484
rect 1276 1476 1284 1484
rect 1292 1476 1300 1484
rect 1548 1476 1556 1484
rect 2060 1476 2068 1484
rect 1212 1456 1220 1464
rect 1100 1416 1108 1424
rect 1164 1416 1172 1424
rect 1516 1436 1524 1444
rect 1548 1436 1556 1444
rect 1740 1436 1748 1444
rect 1788 1436 1796 1444
rect 1694 1406 1702 1414
rect 1708 1406 1716 1414
rect 1722 1406 1730 1414
rect 1276 1336 1284 1344
rect 1324 1336 1332 1344
rect 1516 1336 1524 1344
rect 780 1316 788 1324
rect 828 1316 836 1324
rect 748 1096 756 1104
rect 748 1076 756 1084
rect 748 1056 756 1064
rect 732 1036 740 1044
rect 764 1036 772 1044
rect 748 976 756 984
rect 748 956 756 964
rect 668 916 676 924
rect 940 1236 948 1244
rect 1020 1256 1028 1264
rect 1132 1316 1140 1324
rect 1196 1316 1204 1324
rect 1068 1256 1076 1264
rect 1052 1176 1060 1184
rect 988 1156 996 1164
rect 1036 1156 1044 1164
rect 908 1136 916 1144
rect 972 1136 980 1144
rect 812 1116 820 1124
rect 796 1036 804 1044
rect 940 1116 948 1124
rect 1020 1116 1028 1124
rect 892 1096 900 1104
rect 956 1096 964 1104
rect 1052 1116 1060 1124
rect 892 1076 900 1084
rect 860 1056 868 1064
rect 908 1036 916 1044
rect 828 1016 836 1024
rect 796 996 804 1004
rect 844 996 852 1004
rect 460 876 468 884
rect 668 836 676 844
rect 686 806 694 814
rect 700 806 708 814
rect 714 806 722 814
rect 12 696 20 704
rect 364 696 372 704
rect 476 696 484 704
rect 508 696 516 704
rect 236 656 244 664
rect 28 556 36 564
rect 60 556 68 564
rect 12 496 20 504
rect 268 616 276 624
rect 316 616 324 624
rect 252 596 260 604
rect 188 576 196 584
rect 300 576 308 584
rect 108 556 116 564
rect 124 556 132 564
rect 204 556 212 564
rect 252 556 260 564
rect 92 536 100 544
rect 140 536 148 544
rect 268 536 276 544
rect 364 536 372 544
rect 236 516 244 524
rect 380 516 388 524
rect 396 516 404 524
rect 428 516 436 524
rect 76 496 84 504
rect 364 496 372 504
rect 316 296 324 304
rect 188 256 196 264
rect 28 176 36 184
rect 364 176 372 184
rect 220 116 228 124
rect 588 656 596 664
rect 588 556 596 564
rect 652 556 660 564
rect 780 916 788 924
rect 860 976 868 984
rect 812 916 820 924
rect 780 876 788 884
rect 796 836 804 844
rect 492 536 500 544
rect 556 536 564 544
rect 748 536 756 544
rect 892 956 900 964
rect 988 996 996 1004
rect 956 916 964 924
rect 988 916 996 924
rect 1020 956 1028 964
rect 1004 876 1012 884
rect 876 836 884 844
rect 1084 1156 1092 1164
rect 1196 1296 1204 1304
rect 1292 1296 1300 1304
rect 1148 1136 1156 1144
rect 1164 1136 1172 1144
rect 1100 1056 1108 1064
rect 1100 1016 1108 1024
rect 1084 996 1092 1004
rect 1084 956 1092 964
rect 972 656 980 664
rect 940 636 948 644
rect 1180 1076 1188 1084
rect 1132 996 1140 1004
rect 1180 996 1188 1004
rect 1132 956 1140 964
rect 1164 956 1172 964
rect 1292 1276 1300 1284
rect 1244 1156 1252 1164
rect 1276 1136 1284 1144
rect 1372 1256 1380 1264
rect 1420 1256 1428 1264
rect 1340 1136 1348 1144
rect 1292 1116 1300 1124
rect 1324 1116 1332 1124
rect 1244 1096 1252 1104
rect 1292 1056 1300 1064
rect 1244 1016 1252 1024
rect 1324 1036 1332 1044
rect 1308 1016 1316 1024
rect 1772 1336 1780 1344
rect 2204 1776 2212 1784
rect 2380 1776 2388 1784
rect 2348 1756 2356 1764
rect 2204 1736 2212 1744
rect 2236 1736 2244 1744
rect 2284 1736 2292 1744
rect 2284 1716 2292 1724
rect 2332 1716 2340 1724
rect 2252 1576 2260 1584
rect 2204 1476 2212 1484
rect 2252 1456 2260 1464
rect 2284 1576 2292 1584
rect 2348 1576 2356 1584
rect 2300 1496 2308 1504
rect 2332 1496 2340 1504
rect 2028 1436 2036 1444
rect 2188 1436 2196 1444
rect 1980 1376 1988 1384
rect 2156 1376 2164 1384
rect 1820 1316 1828 1324
rect 1708 1296 1716 1304
rect 1900 1336 1908 1344
rect 2012 1336 2020 1344
rect 2332 1336 2340 1344
rect 2348 1336 2350 1344
rect 2350 1336 2356 1344
rect 1916 1316 1924 1324
rect 1852 1296 1860 1304
rect 1788 1276 1796 1284
rect 1484 1216 1492 1224
rect 1548 1216 1556 1224
rect 1644 1136 1652 1144
rect 1820 1136 1828 1144
rect 1756 1116 1764 1124
rect 1452 1056 1460 1064
rect 1564 1056 1572 1064
rect 1100 936 1108 944
rect 1132 936 1140 944
rect 1228 936 1236 944
rect 1100 916 1108 924
rect 1116 896 1124 904
rect 1180 896 1188 904
rect 1260 896 1268 904
rect 1452 936 1460 944
rect 1436 916 1444 924
rect 1292 856 1300 864
rect 1644 996 1652 1004
rect 1484 976 1492 984
rect 1532 976 1540 984
rect 1580 956 1588 964
rect 1532 936 1540 944
rect 1694 1006 1702 1014
rect 1708 1006 1716 1014
rect 1722 1006 1730 1014
rect 1724 976 1732 984
rect 1740 956 1748 964
rect 1660 936 1668 944
rect 1628 916 1636 924
rect 1644 916 1652 924
rect 1420 836 1428 844
rect 1132 776 1140 784
rect 1196 776 1204 784
rect 1244 776 1252 784
rect 1292 776 1300 784
rect 1116 676 1124 684
rect 1276 676 1284 684
rect 956 616 964 624
rect 1084 616 1092 624
rect 1564 896 1572 904
rect 1596 896 1604 904
rect 1740 916 1748 924
rect 1644 896 1652 904
rect 1596 876 1604 884
rect 1628 876 1636 884
rect 1580 856 1588 864
rect 1532 836 1540 844
rect 1628 836 1636 844
rect 1660 876 1668 884
rect 1724 876 1732 884
rect 1644 736 1652 744
rect 1484 676 1492 684
rect 1148 636 1156 644
rect 844 556 852 564
rect 972 556 980 564
rect 1004 556 1012 564
rect 1036 556 1044 564
rect 1132 556 1140 564
rect 1196 556 1204 564
rect 1244 556 1252 564
rect 876 536 884 544
rect 588 516 596 524
rect 540 476 548 484
rect 604 476 612 484
rect 476 296 484 304
rect 540 296 548 304
rect 686 406 694 414
rect 700 406 708 414
rect 714 406 722 414
rect 748 296 756 304
rect 572 276 580 284
rect 572 256 580 264
rect 732 256 740 264
rect 620 196 628 204
rect 652 196 660 204
rect 412 176 420 184
rect 460 176 468 184
rect 508 136 516 144
rect 924 516 932 524
rect 860 496 868 504
rect 908 496 916 504
rect 1100 536 1108 544
rect 1180 540 1188 544
rect 1180 536 1188 540
rect 1004 516 1012 524
rect 1068 516 1076 524
rect 1100 516 1108 524
rect 1052 496 1060 504
rect 796 196 804 204
rect 892 176 900 184
rect 924 176 932 184
rect 956 176 964 184
rect 812 156 820 164
rect 1036 256 1044 264
rect 1116 296 1124 304
rect 1180 296 1188 304
rect 1068 276 1076 284
rect 1132 280 1140 284
rect 1132 276 1140 280
rect 1068 256 1076 264
rect 1132 176 1140 184
rect 924 156 932 164
rect 1020 156 1028 164
rect 892 136 900 144
rect 972 136 980 144
rect 1100 136 1108 144
rect 1164 136 1172 144
rect 412 116 420 124
rect 700 116 708 124
rect 1052 116 1060 124
rect 1324 536 1332 544
rect 1212 496 1220 504
rect 1212 276 1220 284
rect 1244 176 1252 184
rect 1292 276 1298 284
rect 1298 276 1300 284
rect 1276 256 1284 264
rect 1468 536 1476 544
rect 2252 1176 2260 1184
rect 2268 1136 2276 1144
rect 2300 1136 2308 1144
rect 1884 1096 1892 1104
rect 1772 1076 1780 1084
rect 1788 956 1796 964
rect 1804 956 1812 964
rect 1836 916 1844 924
rect 1756 856 1764 864
rect 1900 1056 1908 1064
rect 1900 1036 1908 1044
rect 2028 1056 2036 1064
rect 1964 1016 1972 1024
rect 1996 1016 2004 1024
rect 2140 1056 2148 1064
rect 2028 996 2036 1004
rect 2108 996 2116 1004
rect 1900 936 1908 944
rect 1868 916 1876 924
rect 2188 1036 2196 1044
rect 2108 956 2116 964
rect 1932 916 1940 924
rect 1916 876 1924 884
rect 1804 836 1812 844
rect 1852 836 1860 844
rect 1852 816 1860 824
rect 1804 736 1812 744
rect 1676 716 1684 724
rect 1964 716 1972 724
rect 1788 696 1796 704
rect 1772 676 1780 684
rect 1820 676 1828 684
rect 1884 676 1892 684
rect 1964 676 1972 684
rect 2108 676 2116 684
rect 2300 836 2308 844
rect 2348 1096 2356 1104
rect 2396 1536 2404 1544
rect 2396 1216 2404 1224
rect 2396 896 2404 904
rect 2300 696 2302 704
rect 2302 696 2308 704
rect 2396 696 2404 704
rect 1692 656 1700 664
rect 1788 656 1796 664
rect 1852 656 1860 664
rect 1932 656 1940 664
rect 1694 606 1702 614
rect 1708 606 1716 614
rect 1722 606 1730 614
rect 1612 536 1620 544
rect 1676 536 1684 544
rect 1740 536 1748 544
rect 1484 276 1492 284
rect 1452 256 1460 264
rect 1484 196 1492 204
rect 1836 496 1844 504
rect 1868 636 1876 644
rect 2140 616 2148 624
rect 2172 616 2180 624
rect 1980 556 1988 564
rect 2140 556 2148 564
rect 1900 496 1908 504
rect 1932 496 1940 504
rect 1964 496 1972 504
rect 1884 456 1892 464
rect 1948 456 1956 464
rect 1996 456 2004 464
rect 2172 536 2180 544
rect 2012 416 2020 424
rect 1868 336 1876 344
rect 2012 316 2020 324
rect 1852 276 1860 284
rect 1788 256 1796 264
rect 1980 256 1988 264
rect 1694 206 1702 214
rect 1708 206 1716 214
rect 1722 206 1730 214
rect 1356 176 1364 184
rect 1820 176 1828 184
rect 1260 136 1268 144
rect 1420 116 1428 124
rect 1820 156 1828 164
rect 1788 136 1796 144
rect 1900 136 1908 144
rect 2060 436 2068 444
rect 2332 436 2340 444
rect 2044 296 2052 304
rect 2108 416 2116 424
rect 2124 336 2132 344
rect 2172 336 2180 344
rect 2220 336 2228 344
rect 2108 296 2116 304
rect 2156 296 2164 304
rect 2268 316 2276 324
rect 2332 316 2340 324
rect 2060 276 2068 284
rect 2204 276 2212 284
rect 2252 276 2260 284
rect 2316 296 2324 304
rect 2236 256 2244 264
rect 2284 256 2292 264
rect 2172 216 2180 224
rect 2140 196 2148 204
rect 2188 196 2196 204
rect 2172 156 2180 164
rect 1580 116 1588 124
rect 1692 116 1700 124
rect 1900 116 1908 124
rect 2028 116 2036 124
rect 2044 116 2052 124
rect 1500 36 1508 44
rect 1532 36 1540 44
rect 924 16 932 24
rect 956 16 964 24
rect 686 6 694 14
rect 700 6 708 14
rect 714 6 722 14
rect 1836 16 1844 24
<< metal3 >>
rect 680 2014 728 2016
rect 680 2006 684 2014
rect 694 2006 700 2014
rect 708 2006 714 2014
rect 724 2006 728 2014
rect 680 2004 728 2006
rect 788 1937 972 1943
rect 980 1937 1084 1943
rect 1028 1917 1228 1923
rect 1396 1917 1564 1923
rect 1892 1917 1932 1923
rect 980 1897 1004 1903
rect 1012 1897 1164 1903
rect 1428 1897 1884 1903
rect 1940 1897 1980 1903
rect 1988 1897 2012 1903
rect 84 1877 220 1883
rect 324 1877 364 1883
rect 372 1877 492 1883
rect 708 1877 1196 1883
rect 1204 1877 1372 1883
rect 1444 1877 1468 1883
rect 1956 1877 2060 1883
rect 820 1857 1148 1863
rect 1156 1857 1260 1863
rect 1300 1857 1596 1863
rect 1604 1857 1852 1863
rect 596 1837 1020 1843
rect 1092 1837 1212 1843
rect 1860 1837 2188 1843
rect 1108 1817 1324 1823
rect 1412 1817 1516 1823
rect 1688 1814 1736 1816
rect 1688 1806 1692 1814
rect 1702 1806 1708 1814
rect 1716 1806 1722 1814
rect 1732 1806 1736 1814
rect 1688 1804 1736 1806
rect 420 1797 444 1803
rect 452 1797 716 1803
rect 724 1797 908 1803
rect 1828 1797 2076 1803
rect 36 1777 380 1783
rect 388 1777 588 1783
rect 596 1777 748 1783
rect 756 1777 924 1783
rect 1588 1777 1932 1783
rect 1972 1777 2204 1783
rect 2212 1777 2380 1783
rect 196 1757 284 1763
rect 772 1757 796 1763
rect 1540 1757 1596 1763
rect 1604 1757 1756 1763
rect 1940 1757 2156 1763
rect 2164 1757 2348 1763
rect 116 1737 652 1743
rect 820 1737 860 1743
rect 868 1737 892 1743
rect 1076 1737 1324 1743
rect 2212 1737 2236 1743
rect 2244 1737 2284 1743
rect 260 1717 460 1723
rect 660 1717 764 1723
rect 1556 1717 1580 1723
rect 2292 1717 2332 1723
rect 772 1697 780 1703
rect 932 1697 1116 1703
rect 1444 1697 1724 1703
rect 1108 1677 1292 1683
rect 1364 1617 1468 1623
rect 680 1614 728 1616
rect 680 1606 684 1614
rect 694 1606 700 1614
rect 708 1606 714 1614
rect 724 1606 728 1614
rect 680 1604 728 1606
rect 724 1577 876 1583
rect 1684 1577 1868 1583
rect 1876 1577 2252 1583
rect 2260 1577 2284 1583
rect 2292 1577 2348 1583
rect 676 1537 828 1543
rect 2404 1537 2435 1543
rect 500 1517 844 1523
rect 1108 1517 1548 1523
rect 324 1497 364 1503
rect 372 1497 380 1503
rect 644 1497 796 1503
rect 804 1497 940 1503
rect 948 1497 972 1503
rect 996 1497 1324 1503
rect 1860 1497 2300 1503
rect 2340 1497 2435 1503
rect 788 1477 812 1483
rect 948 1477 1132 1483
rect 1236 1477 1276 1483
rect 1300 1477 1548 1483
rect 2068 1477 2204 1483
rect 1220 1457 2252 1463
rect 852 1437 908 1443
rect 1524 1437 1548 1443
rect 1748 1437 1788 1443
rect 2036 1437 2188 1443
rect 196 1417 236 1423
rect 244 1417 524 1423
rect 532 1417 620 1423
rect 1108 1417 1164 1423
rect 1688 1414 1736 1416
rect 1688 1406 1692 1414
rect 1702 1406 1708 1414
rect 1716 1406 1722 1414
rect 1732 1406 1736 1414
rect 1688 1404 1736 1406
rect 228 1397 444 1403
rect 756 1377 860 1383
rect 868 1377 956 1383
rect 1988 1377 2156 1383
rect 276 1337 396 1343
rect 420 1337 588 1343
rect 836 1337 876 1343
rect 1284 1337 1324 1343
rect 1524 1337 1772 1343
rect 1908 1337 2012 1343
rect 2020 1337 2332 1343
rect 2340 1337 2348 1343
rect 413 1323 419 1336
rect 52 1317 419 1323
rect 653 1323 659 1336
rect 532 1317 780 1323
rect 788 1317 828 1323
rect 1140 1317 1196 1323
rect 1828 1317 1916 1323
rect -19 1297 12 1303
rect 612 1297 652 1303
rect 660 1297 716 1303
rect 1204 1297 1292 1303
rect 1716 1297 1852 1303
rect 564 1277 652 1283
rect 1300 1277 1788 1283
rect 1028 1257 1068 1263
rect 1076 1257 1372 1263
rect 1380 1257 1420 1263
rect 676 1237 940 1243
rect 1492 1217 1548 1223
rect 2404 1217 2435 1223
rect 680 1214 728 1216
rect 680 1206 684 1214
rect 694 1206 700 1214
rect 708 1206 714 1214
rect 724 1206 728 1214
rect 680 1204 728 1206
rect 340 1177 1052 1183
rect 1060 1177 1516 1183
rect 2260 1177 2435 1183
rect 676 1157 988 1163
rect 1044 1157 1084 1163
rect 1092 1157 1244 1163
rect 916 1137 972 1143
rect 980 1137 1148 1143
rect 1172 1137 1276 1143
rect 1348 1137 1644 1143
rect 1652 1137 1820 1143
rect 1828 1137 2268 1143
rect 2308 1137 2435 1143
rect 84 1117 412 1123
rect 420 1117 524 1123
rect 820 1117 940 1123
rect 1028 1117 1052 1123
rect 1060 1117 1100 1123
rect 1300 1117 1324 1123
rect 1332 1117 1756 1123
rect -19 1097 12 1103
rect 372 1097 524 1103
rect 612 1097 748 1103
rect 900 1097 956 1103
rect 1252 1097 1884 1103
rect 2356 1097 2435 1103
rect 548 1077 748 1083
rect 756 1077 892 1083
rect 1188 1077 1772 1083
rect 580 1057 748 1063
rect 756 1057 860 1063
rect 1300 1057 1452 1063
rect 1572 1057 1900 1063
rect 2036 1057 2140 1063
rect 276 1037 444 1043
rect 516 1037 732 1043
rect 772 1037 796 1043
rect 804 1037 908 1043
rect 916 1037 1324 1043
rect 1908 1037 2188 1043
rect 180 1017 236 1023
rect 644 1017 828 1023
rect 836 1017 1100 1023
rect 1252 1017 1308 1023
rect 1972 1017 1996 1023
rect 1688 1014 1736 1016
rect 1688 1006 1692 1014
rect 1702 1006 1708 1014
rect 1716 1006 1722 1014
rect 1732 1006 1736 1014
rect 1688 1004 1736 1006
rect 804 997 844 1003
rect 852 997 988 1003
rect 1092 997 1132 1003
rect 1188 997 1644 1003
rect 2036 997 2108 1003
rect 52 977 60 983
rect 68 977 444 983
rect 452 977 556 983
rect 564 977 604 983
rect 756 977 860 983
rect 893 977 1484 983
rect 893 964 899 977
rect 1540 977 1724 983
rect -19 957 60 963
rect 68 957 332 963
rect 500 957 572 963
rect 756 957 892 963
rect 1028 957 1084 963
rect 1140 957 1164 963
rect 1588 957 1740 963
rect 1780 957 1788 963
rect 1812 957 2108 963
rect 356 937 460 943
rect 573 943 579 956
rect 573 937 1091 943
rect 564 917 668 923
rect 788 917 812 923
rect 964 917 988 923
rect 1085 923 1091 937
rect 1108 937 1132 943
rect 1140 937 1228 943
rect 1460 937 1532 943
rect 1668 937 1900 943
rect 1085 917 1100 923
rect 1444 917 1628 923
rect 1652 917 1667 923
rect -19 897 12 903
rect 1124 897 1180 903
rect 1188 897 1260 903
rect 1533 897 1564 903
rect 468 877 780 883
rect 1533 883 1539 897
rect 1604 897 1644 903
rect 1661 903 1667 917
rect 1748 917 1836 923
rect 1876 917 1932 923
rect 1661 897 1772 903
rect 2404 897 2435 903
rect 1012 877 1539 883
rect 1549 877 1596 883
rect 1549 863 1555 877
rect 1636 877 1660 883
rect 1732 877 1916 883
rect 1300 857 1555 863
rect 1588 857 1756 863
rect 676 837 796 843
rect 884 837 1420 843
rect 1540 837 1628 843
rect 1812 837 1852 843
rect 1860 837 2300 843
rect 1421 823 1427 836
rect 1421 817 1852 823
rect 680 814 728 816
rect 680 806 684 814
rect 694 806 700 814
rect 708 806 714 814
rect 724 806 728 814
rect 680 804 728 806
rect 1140 777 1196 783
rect 1252 777 1292 783
rect 1300 777 1388 783
rect 1652 737 1804 743
rect 1684 717 1964 723
rect -19 697 12 703
rect 372 697 476 703
rect 484 697 508 703
rect 1796 697 2300 703
rect 2404 697 2435 703
rect 1108 677 1116 683
rect 1284 677 1484 683
rect 1780 677 1820 683
rect 1828 677 1884 683
rect 1972 677 2108 683
rect 244 657 556 663
rect 564 657 588 663
rect 596 657 972 663
rect 1700 657 1788 663
rect 1860 657 1932 663
rect 948 637 1148 643
rect 1780 637 1868 643
rect 276 617 316 623
rect 964 617 1084 623
rect 2148 617 2172 623
rect 1688 614 1736 616
rect 1688 606 1692 614
rect 1702 606 1708 614
rect 1716 606 1722 614
rect 1732 606 1736 614
rect 1688 604 1736 606
rect 20 597 252 603
rect 196 577 300 583
rect -19 557 12 563
rect 36 557 60 563
rect 68 557 108 563
rect 132 557 204 563
rect 260 557 563 563
rect 557 544 563 557
rect 596 557 652 563
rect 852 557 972 563
rect 1012 557 1036 563
rect 1140 557 1196 563
rect 1204 557 1244 563
rect 1988 557 2140 563
rect 100 537 140 543
rect 148 537 268 543
rect 372 537 492 543
rect 564 537 748 543
rect 756 537 876 543
rect 1108 537 1180 543
rect 1332 537 1468 543
rect 1524 537 1612 543
rect 1620 537 1676 543
rect 1748 537 2156 543
rect 2164 537 2172 543
rect 244 517 380 523
rect 404 517 428 523
rect 436 517 588 523
rect 932 517 1004 523
rect 1012 517 1068 523
rect 1076 517 1100 523
rect -19 497 12 503
rect 84 497 364 503
rect 381 503 387 516
rect 381 497 860 503
rect 868 497 908 503
rect 1060 497 1212 503
rect 1844 497 1900 503
rect 1940 497 1964 503
rect 548 477 604 483
rect 1892 457 1948 463
rect 1956 457 1996 463
rect 2068 437 2332 443
rect 2020 417 2108 423
rect 680 414 728 416
rect 680 406 684 414
rect 694 406 700 414
rect 708 406 714 414
rect 724 406 728 414
rect 680 404 728 406
rect 1876 337 2124 343
rect 2132 337 2172 343
rect 2180 337 2220 343
rect 2020 317 2268 323
rect 2276 317 2332 323
rect 324 297 476 303
rect 548 297 748 303
rect 1124 297 1180 303
rect 2052 297 2108 303
rect 2116 297 2156 303
rect 2324 297 2435 303
rect 532 277 572 283
rect 1076 277 1132 283
rect 1140 277 1212 283
rect 1220 277 1292 283
rect 1437 277 1484 283
rect 196 257 556 263
rect 564 257 572 263
rect 580 257 732 263
rect 1044 257 1068 263
rect 1437 263 1443 277
rect 1860 277 2060 283
rect 2212 277 2252 283
rect 1284 257 1443 263
rect 1460 257 1788 263
rect 1988 257 2236 263
rect 2244 257 2284 263
rect 2164 217 2172 223
rect 1688 214 1736 216
rect 1688 206 1692 214
rect 1702 206 1708 214
rect 1716 206 1722 214
rect 1732 206 1736 214
rect 1688 204 1736 206
rect 628 197 652 203
rect 804 197 1484 203
rect 2148 197 2188 203
rect 36 177 364 183
rect 372 177 412 183
rect 420 177 460 183
rect 900 177 924 183
rect 964 177 1132 183
rect 1140 177 1244 183
rect 1252 177 1356 183
rect 1828 177 1836 183
rect 820 157 924 163
rect 932 157 1020 163
rect 1828 157 2172 163
rect 516 137 524 143
rect 900 137 972 143
rect 980 137 1100 143
rect 1172 137 1260 143
rect 1796 137 1900 143
rect 228 117 412 123
rect 708 117 1052 123
rect 1396 117 1420 123
rect 1588 117 1692 123
rect 1908 117 2028 123
rect 2036 117 2044 123
rect 1508 37 1532 43
rect 932 17 956 23
rect 680 14 728 16
rect 680 6 684 14
rect 694 6 700 14
rect 708 6 714 14
rect 724 6 728 14
rect 680 4 728 6
<< m4contact >>
rect 684 2006 686 2014
rect 686 2006 692 2014
rect 700 2006 708 2014
rect 716 2006 722 2014
rect 722 2006 724 2014
rect 780 1996 788 2004
rect 972 1936 980 1944
rect 1932 1916 1940 1924
rect 1692 1806 1694 1814
rect 1694 1806 1700 1814
rect 1708 1806 1716 1814
rect 1724 1806 1730 1814
rect 1730 1806 1732 1814
rect 1932 1756 1940 1764
rect 972 1736 980 1744
rect 780 1696 788 1704
rect 684 1606 686 1614
rect 686 1606 692 1614
rect 700 1606 708 1614
rect 716 1606 722 1614
rect 722 1606 724 1614
rect 1100 1516 1108 1524
rect 1692 1406 1694 1414
rect 1694 1406 1700 1414
rect 1708 1406 1716 1414
rect 1724 1406 1730 1414
rect 1730 1406 1732 1414
rect 684 1206 686 1214
rect 686 1206 692 1214
rect 700 1206 708 1214
rect 716 1206 722 1214
rect 722 1206 724 1214
rect 1516 1176 1524 1184
rect 1100 1116 1108 1124
rect 1100 1056 1108 1064
rect 1692 1006 1694 1014
rect 1694 1006 1700 1014
rect 1708 1006 1716 1014
rect 1724 1006 1730 1014
rect 1730 1006 1732 1014
rect 1772 956 1780 964
rect 1772 896 1780 904
rect 684 806 686 814
rect 686 806 692 814
rect 700 806 708 814
rect 716 806 722 814
rect 722 806 724 814
rect 1388 776 1396 784
rect 1100 676 1108 684
rect 556 656 564 664
rect 1772 636 1780 644
rect 1692 606 1694 614
rect 1694 606 1700 614
rect 1708 606 1716 614
rect 1724 606 1730 614
rect 1730 606 1732 614
rect 12 596 20 604
rect 12 556 20 564
rect 1516 536 1524 544
rect 2156 536 2164 544
rect 684 406 686 414
rect 686 406 692 414
rect 700 406 708 414
rect 716 406 722 414
rect 722 406 724 414
rect 524 276 532 284
rect 556 256 564 264
rect 2156 216 2164 224
rect 1692 206 1694 214
rect 1694 206 1700 214
rect 1708 206 1716 214
rect 1724 206 1730 214
rect 1730 206 1732 214
rect 1836 176 1844 184
rect 524 136 532 144
rect 1388 116 1396 124
rect 1836 16 1844 24
rect 684 6 686 14
rect 686 6 692 14
rect 700 6 708 14
rect 716 6 722 14
rect 722 6 724 14
<< metal4 >>
rect 680 2014 728 2040
rect 680 2006 684 2014
rect 692 2006 700 2014
rect 708 2006 716 2014
rect 724 2006 728 2014
rect 680 1614 728 2006
rect 778 2004 790 2006
rect 778 1996 780 2004
rect 788 1996 790 2004
rect 778 1704 790 1996
rect 970 1944 982 1946
rect 970 1936 972 1944
rect 980 1936 982 1944
rect 970 1744 982 1936
rect 970 1736 972 1744
rect 980 1736 982 1744
rect 970 1734 982 1736
rect 1688 1814 1736 2040
rect 1688 1806 1692 1814
rect 1700 1806 1708 1814
rect 1716 1806 1724 1814
rect 1732 1806 1736 1814
rect 778 1696 780 1704
rect 788 1696 790 1704
rect 778 1694 790 1696
rect 680 1606 684 1614
rect 692 1606 700 1614
rect 708 1606 716 1614
rect 724 1606 728 1614
rect 680 1214 728 1606
rect 680 1206 684 1214
rect 692 1206 700 1214
rect 708 1206 716 1214
rect 724 1206 728 1214
rect 680 814 728 1206
rect 1098 1524 1110 1526
rect 1098 1516 1100 1524
rect 1108 1516 1110 1524
rect 1098 1124 1110 1516
rect 1688 1414 1736 1806
rect 1930 1924 1942 1926
rect 1930 1916 1932 1924
rect 1940 1916 1942 1924
rect 1930 1764 1942 1916
rect 1930 1756 1932 1764
rect 1940 1756 1942 1764
rect 1930 1754 1942 1756
rect 1688 1406 1692 1414
rect 1700 1406 1708 1414
rect 1716 1406 1724 1414
rect 1732 1406 1736 1414
rect 1098 1116 1100 1124
rect 1108 1116 1110 1124
rect 1098 1114 1110 1116
rect 1514 1184 1526 1186
rect 1514 1176 1516 1184
rect 1524 1176 1526 1184
rect 680 806 684 814
rect 692 806 700 814
rect 708 806 716 814
rect 724 806 728 814
rect 554 664 566 666
rect 554 656 556 664
rect 564 656 566 664
rect 10 604 22 606
rect 10 596 12 604
rect 20 596 22 604
rect 10 564 22 596
rect 10 556 12 564
rect 20 556 22 564
rect 10 554 22 556
rect 522 284 534 286
rect 522 276 524 284
rect 532 276 534 284
rect 522 144 534 276
rect 554 264 566 656
rect 554 256 556 264
rect 564 256 566 264
rect 554 254 566 256
rect 680 414 728 806
rect 1098 1064 1110 1066
rect 1098 1056 1100 1064
rect 1108 1056 1110 1064
rect 1098 684 1110 1056
rect 1098 676 1100 684
rect 1108 676 1110 684
rect 1098 674 1110 676
rect 1386 784 1398 786
rect 1386 776 1388 784
rect 1396 776 1398 784
rect 680 406 684 414
rect 692 406 700 414
rect 708 406 716 414
rect 724 406 728 414
rect 522 136 524 144
rect 532 136 534 144
rect 522 134 534 136
rect 680 14 728 406
rect 1386 124 1398 776
rect 1514 544 1526 1176
rect 1514 536 1516 544
rect 1524 536 1526 544
rect 1514 534 1526 536
rect 1688 1014 1736 1406
rect 1688 1006 1692 1014
rect 1700 1006 1708 1014
rect 1716 1006 1724 1014
rect 1732 1006 1736 1014
rect 1688 614 1736 1006
rect 1770 964 1782 966
rect 1770 956 1772 964
rect 1780 956 1782 964
rect 1770 904 1782 956
rect 1770 896 1772 904
rect 1780 896 1782 904
rect 1770 644 1782 896
rect 1770 636 1772 644
rect 1780 636 1782 644
rect 1770 634 1782 636
rect 1688 606 1692 614
rect 1700 606 1708 614
rect 1716 606 1724 614
rect 1732 606 1736 614
rect 1386 116 1388 124
rect 1396 116 1398 124
rect 1386 114 1398 116
rect 1688 214 1736 606
rect 2154 544 2166 546
rect 2154 536 2156 544
rect 2164 536 2166 544
rect 2154 224 2166 536
rect 2154 216 2156 224
rect 2164 216 2166 224
rect 2154 214 2166 216
rect 1688 206 1692 214
rect 1700 206 1708 214
rect 1716 206 1724 214
rect 1732 206 1736 214
rect 680 6 684 14
rect 692 6 700 14
rect 708 6 716 14
rect 724 6 728 14
rect 680 -40 728 6
rect 1688 -40 1736 206
rect 1834 184 1846 186
rect 1834 176 1836 184
rect 1844 176 1846 184
rect 1834 24 1846 176
rect 1834 16 1836 24
rect 1844 16 1846 24
rect 1834 14 1846 16
use DFFSR  DFFSR_2
timestamp 1745250350
transform -1 0 360 0 -1 210
box -4 -6 356 206
use BUFX2  BUFX2_2
timestamp 1745250350
transform 1 0 360 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_4
timestamp 1745250350
transform -1 0 360 0 1 210
box -4 -6 356 206
use BUFX2  BUFX2_1
timestamp 1745250350
transform -1 0 408 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_1
timestamp 1745250350
transform -1 0 520 0 -1 210
box -4 -6 116 206
use FILL  FILL_0_0_0
timestamp 1745250350
transform 1 0 520 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1745250350
transform 1 0 536 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1745250350
transform 1 0 552 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_8
timestamp 1745250350
transform 1 0 568 0 -1 210
box -4 -6 356 206
use DFFSR  DFFSR_5
timestamp 1745250350
transform 1 0 408 0 1 210
box -4 -6 356 206
use XNOR2X1  XNOR2X1_3
timestamp 1745250350
transform -1 0 920 0 1 210
box -4 -6 116 206
use FILL  FILL_1_0_2
timestamp 1745250350
transform -1 0 808 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1745250350
transform -1 0 792 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_0
timestamp 1745250350
transform -1 0 776 0 1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_2
timestamp 1745250350
transform -1 0 1016 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_4
timestamp 1745250350
transform 1 0 920 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1745250350
transform 1 0 968 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_5
timestamp 1745250350
transform 1 0 920 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_12
timestamp 1745250350
transform 1 0 1064 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_3
timestamp 1745250350
transform -1 0 1064 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_16
timestamp 1745250350
transform 1 0 1048 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_6
timestamp 1745250350
transform 1 0 1016 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_14
timestamp 1745250350
transform 1 0 1224 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_13
timestamp 1745250350
transform -1 0 1224 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_3
timestamp 1745250350
transform 1 0 1112 0 1 210
box -4 -6 68 206
use XOR2X1  XOR2X1_1
timestamp 1745250350
transform 1 0 1256 0 -1 210
box -4 -6 116 206
use BUFX2  BUFX2_6
timestamp 1745250350
transform 1 0 1208 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_9
timestamp 1745250350
transform -1 0 1208 0 -1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_3
timestamp 1745250350
transform -1 0 1160 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_10
timestamp 1745250350
transform 1 0 1416 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_7
timestamp 1745250350
transform 1 0 1368 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_6
timestamp 1745250350
transform -1 0 1624 0 1 210
box -4 -6 356 206
use FILL  FILL_1_1_0
timestamp 1745250350
transform 1 0 1624 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1745250350
transform 1 0 1624 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1745250350
transform 1 0 1608 0 -1 210
box -4 -6 20 206
use BUFX4  BUFX4_5
timestamp 1745250350
transform 1 0 1544 0 -1 210
box -4 -6 68 206
use INVX8  INVX8_1
timestamp 1745250350
transform -1 0 1544 0 -1 210
box -4 -6 84 206
use CLKBUF1  CLKBUF1_5
timestamp 1745250350
transform 1 0 1672 0 1 210
box -4 -6 148 206
use FILL  FILL_1_1_2
timestamp 1745250350
transform 1 0 1656 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1745250350
transform 1 0 1640 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1745250350
transform 1 0 1640 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_28
timestamp 1745250350
transform 1 0 1656 0 -1 210
box -4 -6 356 206
use DFFSR  DFFSR_29
timestamp 1745250350
transform 1 0 2008 0 -1 210
box -4 -6 356 206
use BUFX2  BUFX2_30
timestamp 1745250350
transform -1 0 1864 0 1 210
box -4 -6 52 206
use XOR2X1  XOR2X1_8
timestamp 1745250350
transform 1 0 1864 0 1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_12
timestamp 1745250350
transform 1 0 1976 0 1 210
box -4 -6 52 206
use INVX1  INVX1_20
timestamp 1745250350
transform 1 0 2024 0 1 210
box -4 -6 36 206
use INVX1  INVX1_21
timestamp 1745250350
transform 1 0 2056 0 1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_13
timestamp 1745250350
transform 1 0 2088 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_6
timestamp 1745250350
transform 1 0 2152 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1
timestamp 1745250350
transform -1 0 2376 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_2
timestamp 1745250350
transform -1 0 2392 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_3
timestamp 1745250350
transform -1 0 2408 0 -1 210
box -4 -6 20 206
use AOI21X1  AOI21X1_5
timestamp 1745250350
transform 1 0 2216 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_28
timestamp 1745250350
transform 1 0 2280 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_29
timestamp 1745250350
transform 1 0 2328 0 1 210
box -4 -6 52 206
use FILL  FILL_2_1
timestamp 1745250350
transform 1 0 2376 0 1 210
box -4 -6 20 206
use FILL  FILL_2_2
timestamp 1745250350
transform 1 0 2392 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_4
timestamp 1745250350
transform -1 0 56 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_2
timestamp 1745250350
transform 1 0 56 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_1
timestamp 1745250350
transform -1 0 168 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_5
timestamp 1745250350
transform -1 0 200 0 -1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_2
timestamp 1745250350
transform -1 0 264 0 -1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_2
timestamp 1745250350
transform -1 0 376 0 -1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_1
timestamp 1745250350
transform -1 0 472 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_1
timestamp 1745250350
transform -1 0 424 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_19
timestamp 1745250350
transform 1 0 472 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1745250350
transform -1 0 552 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_18
timestamp 1745250350
transform -1 0 600 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_10
timestamp 1745250350
transform 1 0 648 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_11
timestamp 1745250350
transform -1 0 648 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_0_0
timestamp 1745250350
transform -1 0 712 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1745250350
transform -1 0 744 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1745250350
transform -1 0 728 0 -1 610
box -4 -6 20 206
use BUFX4  BUFX4_4
timestamp 1745250350
transform -1 0 808 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_5
timestamp 1745250350
transform -1 0 872 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_20
timestamp 1745250350
transform 1 0 872 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_5
timestamp 1745250350
transform 1 0 920 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_7
timestamp 1745250350
transform 1 0 968 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_15
timestamp 1745250350
transform -1 0 1048 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_2
timestamp 1745250350
transform 1 0 1048 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1745250350
transform -1 0 1144 0 -1 610
box -4 -6 36 206
use AND2X2  AND2X2_4
timestamp 1745250350
transform -1 0 1208 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1745250350
transform -1 0 1256 0 -1 610
box -4 -6 52 206
use DFFSR  DFFSR_7
timestamp 1745250350
transform -1 0 1608 0 -1 610
box -4 -6 356 206
use CLKBUF1  CLKBUF1_4
timestamp 1745250350
transform 1 0 1608 0 -1 610
box -4 -6 148 206
use FILL  FILL_2_1_0
timestamp 1745250350
transform 1 0 1752 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1745250350
transform 1 0 1768 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1745250350
transform 1 0 1784 0 -1 610
box -4 -6 20 206
use NAND2X1  NAND2X1_13
timestamp 1745250350
transform 1 0 1800 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_7
timestamp 1745250350
transform -1 0 1896 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_5
timestamp 1745250350
transform -1 0 1960 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_30
timestamp 1745250350
transform -1 0 2008 0 -1 610
box -4 -6 52 206
use DFFSR  DFFSR_30
timestamp 1745250350
transform 1 0 2008 0 -1 610
box -4 -6 356 206
use FILL  FILL_3_1
timestamp 1745250350
transform -1 0 2376 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_2
timestamp 1745250350
transform -1 0 2392 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_3
timestamp 1745250350
transform -1 0 2408 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_3
timestamp 1745250350
transform -1 0 56 0 1 610
box -4 -6 52 206
use DFFSR  DFFSR_3
timestamp 1745250350
transform -1 0 408 0 1 610
box -4 -6 356 206
use DFFSR  DFFSR_1
timestamp 1745250350
transform -1 0 760 0 1 610
box -4 -6 356 206
use FILL  FILL_3_0_0
timestamp 1745250350
transform 1 0 760 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1745250350
transform 1 0 776 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1745250350
transform 1 0 792 0 1 610
box -4 -6 20 206
use DFFSR  DFFSR_9
timestamp 1745250350
transform 1 0 808 0 1 610
box -4 -6 356 206
use XNOR2X1  XNOR2X1_4
timestamp 1745250350
transform 1 0 1160 0 1 610
box -4 -6 116 206
use DFFSR  DFFSR_10
timestamp 1745250350
transform -1 0 1624 0 1 610
box -4 -6 356 206
use INVX1  INVX1_19
timestamp 1745250350
transform -1 0 1656 0 1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_32
timestamp 1745250350
transform -1 0 1704 0 1 610
box -4 -6 52 206
use FILL  FILL_3_1_0
timestamp 1745250350
transform -1 0 1720 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1745250350
transform -1 0 1736 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1745250350
transform -1 0 1752 0 1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_12
timestamp 1745250350
transform -1 0 1816 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_33
timestamp 1745250350
transform 1 0 1816 0 1 610
box -4 -6 52 206
use OR2X2  OR2X2_1
timestamp 1745250350
transform 1 0 1864 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_34
timestamp 1745250350
transform 1 0 1928 0 1 610
box -4 -6 52 206
use DFFSR  DFFSR_27
timestamp 1745250350
transform 1 0 1976 0 1 610
box -4 -6 356 206
use BUFX2  BUFX2_12
timestamp 1745250350
transform 1 0 2328 0 1 610
box -4 -6 52 206
use FILL  FILL_4_1
timestamp 1745250350
transform 1 0 2376 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1745250350
transform 1 0 2392 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_24
timestamp 1745250350
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use CLKBUF1  CLKBUF1_2
timestamp 1745250350
transform 1 0 56 0 -1 1010
box -4 -6 148 206
use CLKBUF1  CLKBUF1_1
timestamp 1745250350
transform -1 0 344 0 -1 1010
box -4 -6 148 206
use XOR2X1  XOR2X1_6
timestamp 1745250350
transform 1 0 344 0 -1 1010
box -4 -6 116 206
use NOR2X1  NOR2X1_30
timestamp 1745250350
transform -1 0 504 0 -1 1010
box -4 -6 52 206
use BUFX4  BUFX4_2
timestamp 1745250350
transform -1 0 568 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_2
timestamp 1745250350
transform -1 0 600 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_8
timestamp 1745250350
transform 1 0 600 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1745250350
transform -1 0 680 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1745250350
transform -1 0 696 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1745250350
transform -1 0 712 0 -1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_31
timestamp 1745250350
transform -1 0 760 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_4
timestamp 1745250350
transform 1 0 760 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_11
timestamp 1745250350
transform 1 0 824 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_17
timestamp 1745250350
transform -1 0 920 0 -1 1010
box -4 -6 36 206
use NOR3X1  NOR3X1_1
timestamp 1745250350
transform -1 0 1048 0 -1 1010
box -4 -6 132 206
use NOR2X1  NOR2X1_5
timestamp 1745250350
transform -1 0 1096 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_9
timestamp 1745250350
transform -1 0 1144 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_17
timestamp 1745250350
transform 1 0 1144 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_6
timestamp 1745250350
transform -1 0 1240 0 -1 1010
box -4 -6 52 206
use AOI22X1  AOI22X1_1
timestamp 1745250350
transform 1 0 1240 0 -1 1010
box -4 -6 84 206
use INVX1  INVX1_24
timestamp 1745250350
transform -1 0 1352 0 -1 1010
box -4 -6 36 206
use NOR3X1  NOR3X1_3
timestamp 1745250350
transform -1 0 1480 0 -1 1010
box -4 -6 132 206
use OAI21X1  OAI21X1_4
timestamp 1745250350
transform 1 0 1480 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1745250350
transform -1 0 1608 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_14
timestamp 1745250350
transform -1 0 1672 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_1_0
timestamp 1745250350
transform 1 0 1672 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1745250350
transform 1 0 1688 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1745250350
transform 1 0 1704 0 -1 1010
box -4 -6 20 206
use AND2X2  AND2X2_7
timestamp 1745250350
transform 1 0 1720 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_23
timestamp 1745250350
transform 1 0 1784 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_6
timestamp 1745250350
transform 1 0 1816 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_22
timestamp 1745250350
transform -1 0 1912 0 -1 1010
box -4 -6 36 206
use AND2X2  AND2X2_8
timestamp 1745250350
transform 1 0 1912 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_26
timestamp 1745250350
transform 1 0 1976 0 -1 1010
box -4 -6 356 206
use BUFX2  BUFX2_27
timestamp 1745250350
transform 1 0 2328 0 -1 1010
box -4 -6 52 206
use FILL  FILL_5_1
timestamp 1745250350
transform -1 0 2392 0 -1 1010
box -4 -6 20 206
use FILL  FILL_5_2
timestamp 1745250350
transform -1 0 2408 0 -1 1010
box -4 -6 20 206
use BUFX2  BUFX2_25
timestamp 1745250350
transform -1 0 56 0 1 1010
box -4 -6 52 206
use DFFSR  DFFSR_25
timestamp 1745250350
transform -1 0 408 0 1 1010
box -4 -6 356 206
use XOR2X1  XOR2X1_7
timestamp 1745250350
transform -1 0 520 0 1 1010
box -4 -6 116 206
use NAND2X1  NAND2X1_14
timestamp 1745250350
transform -1 0 568 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_6
timestamp 1745250350
transform 1 0 568 0 1 1010
box -4 -6 52 206
use FILL  FILL_5_0_0
timestamp 1745250350
transform -1 0 632 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1745250350
transform -1 0 648 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1745250350
transform -1 0 664 0 1 1010
box -4 -6 20 206
use NOR3X1  NOR3X1_2
timestamp 1745250350
transform -1 0 792 0 1 1010
box -4 -6 132 206
use NAND3X1  NAND3X1_6
timestamp 1745250350
transform 1 0 792 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_18
timestamp 1745250350
transform 1 0 856 0 1 1010
box -4 -6 36 206
use INVX1  INVX1_3
timestamp 1745250350
transform 1 0 888 0 1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_9
timestamp 1745250350
transform -1 0 984 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_6
timestamp 1745250350
transform -1 0 1048 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_10
timestamp 1745250350
transform -1 0 1096 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1745250350
transform 1 0 1096 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_2
timestamp 1745250350
transform 1 0 1144 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_3
timestamp 1745250350
transform 1 0 1208 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_3
timestamp 1745250350
transform -1 0 1320 0 1 1010
box -4 -6 68 206
use DFFSR  DFFSR_32
timestamp 1745250350
transform 1 0 1320 0 1 1010
box -4 -6 356 206
use FILL  FILL_5_1_0
timestamp 1745250350
transform 1 0 1672 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1745250350
transform 1 0 1688 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1745250350
transform 1 0 1704 0 1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_15
timestamp 1745250350
transform 1 0 1720 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_8
timestamp 1745250350
transform 1 0 1768 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_16
timestamp 1745250350
transform -1 0 1864 0 1 1010
box -4 -6 52 206
use DFFSR  DFFSR_31
timestamp 1745250350
transform 1 0 1864 0 1 1010
box -4 -6 356 206
use BUFX2  BUFX2_31
timestamp 1745250350
transform 1 0 2216 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_32
timestamp 1745250350
transform 1 0 2264 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_26
timestamp 1745250350
transform 1 0 2312 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_14
timestamp 1745250350
transform 1 0 2360 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_23
timestamp 1745250350
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use DFFSR  DFFSR_24
timestamp 1745250350
transform -1 0 408 0 -1 1410
box -4 -6 356 206
use XOR2X1  XOR2X1_5
timestamp 1745250350
transform -1 0 520 0 -1 1410
box -4 -6 116 206
use NOR2X1  NOR2X1_29
timestamp 1745250350
transform -1 0 568 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_1
timestamp 1745250350
transform -1 0 632 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_7
timestamp 1745250350
transform 1 0 632 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_0_0
timestamp 1745250350
transform 1 0 696 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1745250350
transform 1 0 712 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1745250350
transform 1 0 728 0 -1 1410
box -4 -6 20 206
use INVX1  INVX1_16
timestamp 1745250350
transform 1 0 744 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_28
timestamp 1745250350
transform 1 0 776 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_26
timestamp 1745250350
transform -1 0 872 0 -1 1410
box -4 -6 52 206
use XOR2X1  XOR2X1_4
timestamp 1745250350
transform 1 0 872 0 -1 1410
box -4 -6 116 206
use BUFX4  BUFX4_1
timestamp 1745250350
transform 1 0 984 0 -1 1410
box -4 -6 68 206
use CLKBUF1  CLKBUF1_3
timestamp 1745250350
transform 1 0 1048 0 -1 1410
box -4 -6 148 206
use NOR2X1  NOR2X1_19
timestamp 1745250350
transform -1 0 1240 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_22
timestamp 1745250350
transform -1 0 1288 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1745250350
transform -1 0 1352 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_1
timestamp 1745250350
transform -1 0 1384 0 -1 1410
box -4 -6 36 206
use DFFSR  DFFSR_11
timestamp 1745250350
transform 1 0 1384 0 -1 1410
box -4 -6 356 206
use FILL  FILL_6_1_0
timestamp 1745250350
transform -1 0 1752 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1745250350
transform -1 0 1768 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1745250350
transform -1 0 1784 0 -1 1410
box -4 -6 20 206
use NOR2X1  NOR2X1_18
timestamp 1745250350
transform -1 0 1832 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_9
timestamp 1745250350
transform -1 0 1864 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_7
timestamp 1745250350
transform -1 0 1912 0 -1 1410
box -4 -6 52 206
use XOR2X1  XOR2X1_2
timestamp 1745250350
transform 1 0 1912 0 -1 1410
box -4 -6 116 206
use DFFSR  DFFSR_12
timestamp 1745250350
transform 1 0 2024 0 -1 1410
box -4 -6 356 206
use FILL  FILL_7_1
timestamp 1745250350
transform -1 0 2392 0 -1 1410
box -4 -6 20 206
use FILL  FILL_7_2
timestamp 1745250350
transform -1 0 2408 0 -1 1410
box -4 -6 20 206
use DFFSR  DFFSR_23
timestamp 1745250350
transform -1 0 360 0 1 1410
box -4 -6 356 206
use DFFSR  DFFSR_21
timestamp 1745250350
transform 1 0 360 0 1 1410
box -4 -6 356 206
use FILL  FILL_7_0_0
timestamp 1745250350
transform -1 0 728 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1745250350
transform -1 0 744 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1745250350
transform -1 0 760 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_22
timestamp 1745250350
transform -1 0 808 0 1 1410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_9
timestamp 1745250350
transform -1 0 920 0 1 1410
box -4 -6 116 206
use DFFSR  DFFSR_22
timestamp 1745250350
transform -1 0 1272 0 1 1410
box -4 -6 356 206
use BUFX4  BUFX4_3
timestamp 1745250350
transform -1 0 1336 0 1 1410
box -4 -6 68 206
use DFFSR  DFFSR_33
timestamp 1745250350
transform -1 0 1688 0 1 1410
box -4 -6 356 206
use FILL  FILL_7_1_0
timestamp 1745250350
transform 1 0 1688 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1745250350
transform 1 0 1704 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1745250350
transform 1 0 1720 0 1 1410
box -4 -6 20 206
use XNOR2X1  XNOR2X1_5
timestamp 1745250350
transform 1 0 1736 0 1 1410
box -4 -6 116 206
use DFFSR  DFFSR_13
timestamp 1745250350
transform -1 0 2200 0 1 1410
box -4 -6 356 206
use NOR2X1  NOR2X1_21
timestamp 1745250350
transform -1 0 2248 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_20
timestamp 1745250350
transform -1 0 2296 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_11
timestamp 1745250350
transform 1 0 2296 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_13
timestamp 1745250350
transform 1 0 2344 0 1 1410
box -4 -6 52 206
use FILL  FILL_8_1
timestamp 1745250350
transform 1 0 2392 0 1 1410
box -4 -6 20 206
use XNOR2X1  XNOR2X1_6
timestamp 1745250350
transform -1 0 120 0 -1 1810
box -4 -6 116 206
use DFFSR  DFFSR_18
timestamp 1745250350
transform 1 0 120 0 -1 1810
box -4 -6 356 206
use XNOR2X1  XNOR2X1_7
timestamp 1745250350
transform -1 0 584 0 -1 1810
box -4 -6 116 206
use NAND2X1  NAND2X1_25
timestamp 1745250350
transform 1 0 584 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_13
timestamp 1745250350
transform -1 0 664 0 -1 1810
box -4 -6 36 206
use FILL  FILL_8_0_0
timestamp 1745250350
transform 1 0 664 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1745250350
transform 1 0 680 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1745250350
transform 1 0 696 0 -1 1810
box -4 -6 20 206
use NAND2X1  NAND2X1_26
timestamp 1745250350
transform 1 0 712 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_25
timestamp 1745250350
transform -1 0 808 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_27
timestamp 1745250350
transform 1 0 808 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_29
timestamp 1745250350
transform 1 0 856 0 -1 1810
box -4 -6 52 206
use AND2X2  AND2X2_2
timestamp 1745250350
transform 1 0 904 0 -1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_8
timestamp 1745250350
transform 1 0 968 0 -1 1810
box -4 -6 116 206
use INVX1  INVX1_14
timestamp 1745250350
transform -1 0 1112 0 -1 1810
box -4 -6 36 206
use DFFSR  DFFSR_19
timestamp 1745250350
transform -1 0 1464 0 -1 1810
box -4 -6 356 206
use BUFX2  BUFX2_33
timestamp 1745250350
transform 1 0 1464 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_12
timestamp 1745250350
transform -1 0 1544 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_4
timestamp 1745250350
transform -1 0 1592 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_9
timestamp 1745250350
transform -1 0 1640 0 -1 1810
box -4 -6 52 206
use FILL  FILL_8_1_0
timestamp 1745250350
transform 1 0 1640 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1745250350
transform 1 0 1656 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1745250350
transform 1 0 1672 0 -1 1810
box -4 -6 20 206
use DFFSR  DFFSR_15
timestamp 1745250350
transform 1 0 1688 0 -1 1810
box -4 -6 356 206
use XOR2X1  XOR2X1_3
timestamp 1745250350
transform -1 0 2152 0 -1 1810
box -4 -6 116 206
use NOR2X1  NOR2X1_24
timestamp 1745250350
transform 1 0 2152 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_23
timestamp 1745250350
transform 1 0 2200 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_23
timestamp 1745250350
transform 1 0 2248 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_10
timestamp 1745250350
transform -1 0 2328 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_22
timestamp 1745250350
transform -1 0 2376 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1745250350
transform 1 0 2376 0 -1 1810
box -4 -6 36 206
use DFFSR  DFFSR_17
timestamp 1745250350
transform -1 0 360 0 1 1810
box -4 -6 356 206
use BUFX2  BUFX2_17
timestamp 1745250350
transform 1 0 360 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_18
timestamp 1745250350
transform 1 0 408 0 1 1810
box -4 -6 52 206
use DFFSR  DFFSR_20
timestamp 1745250350
transform 1 0 456 0 1 1810
box -4 -6 356 206
use FILL  FILL_9_0_0
timestamp 1745250350
transform -1 0 824 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1745250350
transform -1 0 840 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1745250350
transform -1 0 856 0 1 1810
box -4 -6 20 206
use BUFX2  BUFX2_21
timestamp 1745250350
transform -1 0 904 0 1 1810
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1745250350
transform 1 0 904 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_11
timestamp 1745250350
transform -1 0 1016 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_28
timestamp 1745250350
transform -1 0 1064 0 1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_5
timestamp 1745250350
transform -1 0 1128 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_15
timestamp 1745250350
transform -1 0 1160 0 1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_27
timestamp 1745250350
transform 1 0 1160 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_3
timestamp 1745250350
transform 1 0 1208 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_20
timestamp 1745250350
transform 1 0 1272 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_19
timestamp 1745250350
transform 1 0 1320 0 1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_4
timestamp 1745250350
transform -1 0 1432 0 1 1810
box -4 -6 68 206
use DFFSR  DFFSR_16
timestamp 1745250350
transform 1 0 1432 0 1 1810
box -4 -6 356 206
use FILL  FILL_9_1_0
timestamp 1745250350
transform 1 0 1784 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1745250350
transform 1 0 1800 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1745250350
transform 1 0 1816 0 1 1810
box -4 -6 20 206
use BUFX2  BUFX2_16
timestamp 1745250350
transform 1 0 1832 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_24
timestamp 1745250350
transform -1 0 1928 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_8
timestamp 1745250350
transform -1 0 1976 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_15
timestamp 1745250350
transform 1 0 1976 0 1 1810
box -4 -6 52 206
use DFFSR  DFFSR_14
timestamp 1745250350
transform 1 0 2024 0 1 1810
box -4 -6 356 206
use FILL  FILL_10_1
timestamp 1745250350
transform 1 0 2376 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_2
timestamp 1745250350
transform 1 0 2392 0 1 1810
box -4 -6 20 206
<< labels >>
flabel metal4 s 680 -40 728 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 1688 -40 1736 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -19 957 -13 963 7 FreeSans 24 0 0 0 clk
port 2 nsew
flabel metal2 s 1501 -23 1507 -17 7 FreeSans 24 270 0 0 reset
port 3 nsew
flabel metal3 s -19 557 -13 563 7 FreeSans 24 0 0 0 enable
port 4 nsew
flabel metal2 s 381 -23 387 -17 7 FreeSans 24 270 0 0 count[0]
port 5 nsew
flabel metal2 s 413 -23 419 -17 7 FreeSans 24 270 0 0 count[1]
port 6 nsew
flabel metal3 s -19 697 -13 703 7 FreeSans 24 0 0 0 count[2]
port 7 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 count[3]
port 8 nsew
flabel metal2 s 925 -23 931 -17 7 FreeSans 24 270 0 0 count[4]
port 9 nsew
flabel metal2 s 1229 -23 1235 -17 7 FreeSans 24 270 0 0 count[5]
port 10 nsew
flabel metal2 s 1389 -23 1395 -17 7 FreeSans 24 270 0 0 count[6]
port 11 nsew
flabel metal2 s 989 -23 995 -17 7 FreeSans 24 270 0 0 count[7]
port 12 nsew
flabel metal2 s 1181 -23 1187 -17 7 FreeSans 24 270 0 0 count[8]
port 13 nsew
flabel metal2 s 1437 -23 1443 -17 7 FreeSans 24 270 0 0 count[9]
port 14 nsew
flabel metal3 s 2429 1497 2435 1503 3 FreeSans 24 0 0 0 count[10]
port 15 nsew
flabel metal3 s 2429 697 2435 703 3 FreeSans 24 0 0 0 count[11]
port 16 nsew
flabel metal3 s 2429 1537 2435 1543 3 FreeSans 24 0 0 0 count[12]
port 17 nsew
flabel metal3 s 2429 1217 2435 1223 3 FreeSans 24 0 0 0 count[13]
port 18 nsew
flabel metal2 s 1997 2037 2003 2043 3 FreeSans 24 90 0 0 count[14]
port 19 nsew
flabel metal2 s 1853 2037 1859 2043 3 FreeSans 24 90 0 0 count[15]
port 20 nsew
flabel metal2 s 381 2037 387 2043 3 FreeSans 24 90 0 0 count[16]
port 21 nsew
flabel metal2 s 429 2037 435 2043 3 FreeSans 24 90 0 0 count[17]
port 22 nsew
flabel metal2 s 1341 2037 1347 2043 3 FreeSans 24 90 0 0 count[18]
port 23 nsew
flabel metal2 s 1293 2037 1299 2043 3 FreeSans 24 90 0 0 count[19]
port 24 nsew
flabel metal2 s 877 2037 883 2043 3 FreeSans 24 90 0 0 count[20]
port 25 nsew
flabel metal2 s 781 2037 787 2043 3 FreeSans 24 90 0 0 count[21]
port 26 nsew
flabel metal3 s -19 1297 -13 1303 7 FreeSans 24 0 0 0 count[22]
port 27 nsew
flabel metal3 s -19 897 -13 903 7 FreeSans 24 0 0 0 count[23]
port 28 nsew
flabel metal3 s -19 1097 -13 1103 7 FreeSans 24 0 0 0 count[24]
port 29 nsew
flabel metal3 s 2429 1097 2435 1103 3 FreeSans 24 0 0 0 count[25]
port 30 nsew
flabel metal3 s 2429 897 2435 903 3 FreeSans 24 0 0 0 count[26]
port 31 nsew
flabel metal3 s 2429 297 2435 303 3 FreeSans 24 0 0 0 count[27]
port 32 nsew
flabel metal2 s 2349 -23 2355 -17 7 FreeSans 24 270 0 0 count[28]
port 33 nsew
flabel metal2 s 1837 -23 1843 -17 7 FreeSans 24 270 0 0 count[29]
port 34 nsew
flabel metal3 s 2429 1177 2435 1183 3 FreeSans 24 0 0 0 count[30]
port 35 nsew
flabel metal3 s 2429 1137 2435 1143 3 FreeSans 24 0 0 0 count[31]
port 36 nsew
flabel metal2 s 1485 2037 1491 2043 3 FreeSans 24 90 0 0 overflow
port 37 nsew
<< end >>
